magic
tech sky130A
magscale 1 2
timestamp 1727525581
<< viali >>
rect 5917 12937 5951 12971
rect 6561 12869 6595 12903
rect 5825 12801 5859 12835
rect 6929 12801 6963 12835
rect 7205 12801 7239 12835
rect 7849 12801 7883 12835
rect 8677 12801 8711 12835
rect 7389 12597 7423 12631
rect 8033 12597 8067 12631
rect 8493 12597 8527 12631
rect 10333 12325 10367 12359
rect 3617 12257 3651 12291
rect 6377 12257 6411 12291
rect 6653 12257 6687 12291
rect 7297 12257 7331 12291
rect 6285 12189 6319 12223
rect 7389 12189 7423 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 10241 12189 10275 12223
rect 10517 12189 10551 12223
rect 10701 12189 10735 12223
rect 1593 12121 1627 12155
rect 3341 12121 3375 12155
rect 5365 12121 5399 12155
rect 9873 12121 9907 12155
rect 10057 12121 10091 12155
rect 5273 12053 5307 12087
rect 7757 12053 7791 12087
rect 7941 12053 7975 12087
rect 2421 11849 2455 11883
rect 4353 11849 4387 11883
rect 8677 11849 8711 11883
rect 9321 11849 9355 11883
rect 9873 11849 9907 11883
rect 2329 11713 2363 11747
rect 2605 11713 2639 11747
rect 4721 11713 4755 11747
rect 4997 11713 5031 11747
rect 5181 11713 5215 11747
rect 5641 11713 5675 11747
rect 5825 11713 5859 11747
rect 5917 11713 5951 11747
rect 8217 11713 8251 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 9505 11713 9539 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10149 11713 10183 11747
rect 10333 11713 10367 11747
rect 10609 11713 10643 11747
rect 10793 11713 10827 11747
rect 11069 11713 11103 11747
rect 2881 11645 2915 11679
rect 4537 11645 4571 11679
rect 5457 11645 5491 11679
rect 5733 11645 5767 11679
rect 7297 11645 7331 11679
rect 7389 11645 7423 11679
rect 7481 11645 7515 11679
rect 7573 11645 7607 11679
rect 8125 11645 8159 11679
rect 8861 11645 8895 11679
rect 9689 11645 9723 11679
rect 7849 11577 7883 11611
rect 10149 11577 10183 11611
rect 7757 11509 7791 11543
rect 8217 11509 8251 11543
rect 3249 11305 3283 11339
rect 4537 11305 4571 11339
rect 4905 11305 4939 11339
rect 7665 11305 7699 11339
rect 7757 11305 7791 11339
rect 10425 11305 10459 11339
rect 11253 11305 11287 11339
rect 1593 11237 1627 11271
rect 10057 11237 10091 11271
rect 4997 11169 5031 11203
rect 5273 11169 5307 11203
rect 7573 11169 7607 11203
rect 10333 11169 10367 11203
rect 10517 11169 10551 11203
rect 11529 11169 11563 11203
rect 11621 11169 11655 11203
rect 1409 11101 1443 11135
rect 3157 11101 3191 11135
rect 4721 11101 4755 11135
rect 5089 11101 5123 11135
rect 5181 11101 5215 11135
rect 5457 11101 5491 11135
rect 5733 11101 5767 11135
rect 5917 11101 5951 11135
rect 7849 11101 7883 11135
rect 10425 11101 10459 11135
rect 10793 11101 10827 11135
rect 10885 11101 10919 11135
rect 10977 11101 11011 11135
rect 11161 11101 11195 11135
rect 11437 11101 11471 11135
rect 11713 11101 11747 11135
rect 5825 11033 5859 11067
rect 5365 10965 5399 10999
rect 6377 10761 6411 10795
rect 10977 10761 11011 10795
rect 1685 10693 1719 10727
rect 3341 10693 3375 10727
rect 8493 10693 8527 10727
rect 8677 10693 8711 10727
rect 10609 10693 10643 10727
rect 11253 10693 11287 10727
rect 3433 10625 3467 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 6561 10625 6595 10659
rect 8125 10625 8159 10659
rect 8217 10625 8251 10659
rect 8401 10625 8435 10659
rect 8861 10625 8895 10659
rect 10793 10625 10827 10659
rect 11069 10625 11103 10659
rect 11345 10625 11379 10659
rect 1409 10557 1443 10591
rect 3157 10557 3191 10591
rect 5089 10557 5123 10591
rect 5549 10557 5583 10591
rect 6837 10557 6871 10591
rect 10701 10557 10735 10591
rect 6009 10489 6043 10523
rect 6745 10489 6779 10523
rect 7941 10489 7975 10523
rect 8309 10421 8343 10455
rect 1501 10217 1535 10251
rect 4997 10217 5031 10251
rect 5549 10217 5583 10251
rect 10149 10217 10183 10251
rect 9413 10149 9447 10183
rect 11805 10149 11839 10183
rect 6101 10081 6135 10115
rect 9873 10081 9907 10115
rect 1685 10013 1719 10047
rect 5181 10013 5215 10047
rect 5365 10013 5399 10047
rect 5457 10013 5491 10047
rect 5733 10013 5767 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 8217 10013 8251 10047
rect 8401 10013 8435 10047
rect 11989 10013 12023 10047
rect 5917 9945 5951 9979
rect 9413 9945 9447 9979
rect 9965 9945 9999 9979
rect 8309 9877 8343 9911
rect 7297 9605 7331 9639
rect 9229 9605 9263 9639
rect 9321 9605 9355 9639
rect 4997 9537 5031 9571
rect 7021 9537 7055 9571
rect 9597 9537 9631 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3249 9469 3283 9503
rect 7297 9469 7331 9503
rect 9689 9469 9723 9503
rect 9873 9401 9907 9435
rect 3157 9333 3191 9367
rect 7113 9333 7147 9367
rect 2421 9129 2455 9163
rect 2881 9129 2915 9163
rect 5917 9129 5951 9163
rect 9137 9129 9171 9163
rect 11897 9129 11931 9163
rect 7757 9061 7791 9095
rect 11161 9061 11195 9095
rect 3249 8993 3283 9027
rect 5733 8993 5767 9027
rect 8309 8993 8343 9027
rect 10057 8993 10091 9027
rect 2605 8925 2639 8959
rect 2973 8925 3007 8959
rect 5641 8925 5675 8959
rect 8953 8925 8987 8959
rect 10149 8925 10183 8959
rect 10977 8925 11011 8959
rect 11161 8925 11195 8959
rect 11805 8925 11839 8959
rect 11989 8925 12023 8959
rect 7481 8857 7515 8891
rect 8125 8857 8159 8891
rect 11345 8857 11379 8891
rect 11529 8857 11563 8891
rect 11713 8857 11747 8891
rect 7573 8789 7607 8823
rect 8217 8789 8251 8823
rect 10517 8789 10551 8823
rect 6009 8585 6043 8619
rect 6377 8585 6411 8619
rect 6929 8585 6963 8619
rect 9229 8585 9263 8619
rect 11897 8585 11931 8619
rect 5365 8517 5399 8551
rect 3341 8449 3375 8483
rect 4813 8449 4847 8483
rect 4997 8449 5031 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 5917 8449 5951 8483
rect 6101 8449 6135 8483
rect 6745 8449 6779 8483
rect 6837 8449 6871 8483
rect 7113 8449 7147 8483
rect 8861 8449 8895 8483
rect 8953 8449 8987 8483
rect 11713 8449 11747 8483
rect 3065 8381 3099 8415
rect 6653 8381 6687 8415
rect 8769 8381 8803 8415
rect 9045 8381 9079 8415
rect 4905 8313 4939 8347
rect 5825 8313 5859 8347
rect 7113 8313 7147 8347
rect 1593 8245 1627 8279
rect 4629 8245 4663 8279
rect 5365 8245 5399 8279
rect 6653 8245 6687 8279
rect 1501 8041 1535 8075
rect 3157 8041 3191 8075
rect 5549 8041 5583 8075
rect 6837 8041 6871 8075
rect 10425 8041 10459 8075
rect 3893 7973 3927 8007
rect 8217 7973 8251 8007
rect 1685 7837 1719 7871
rect 2421 7837 2455 7871
rect 3065 7837 3099 7871
rect 3341 7837 3375 7871
rect 3617 7837 3651 7871
rect 3801 7837 3835 7871
rect 4261 7837 4295 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 10333 7837 10367 7871
rect 10517 7837 10551 7871
rect 6469 7769 6503 7803
rect 8401 7769 8435 7803
rect 3525 7701 3559 7735
rect 6561 7701 6595 7735
rect 6653 7497 6687 7531
rect 7481 7497 7515 7531
rect 9137 7497 9171 7531
rect 10333 7497 10367 7531
rect 7021 7429 7055 7463
rect 8953 7429 8987 7463
rect 3893 7361 3927 7395
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 5089 7361 5123 7395
rect 5457 7361 5491 7395
rect 5641 7361 5675 7395
rect 5733 7361 5767 7395
rect 6193 7361 6227 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 7113 7361 7147 7395
rect 7297 7361 7331 7395
rect 8309 7361 8343 7395
rect 8401 7361 8435 7395
rect 8493 7361 8527 7395
rect 8677 7361 8711 7395
rect 8769 7361 8803 7395
rect 9413 7361 9447 7395
rect 9597 7361 9631 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 10701 7361 10735 7395
rect 10793 7361 10827 7395
rect 10977 7361 11011 7395
rect 4077 7293 4111 7327
rect 3985 7225 4019 7259
rect 9229 7225 9263 7259
rect 3709 7157 3743 7191
rect 6193 7157 6227 7191
rect 8033 7157 8067 7191
rect 9597 7157 9631 7191
rect 6653 6953 6687 6987
rect 9137 6953 9171 6987
rect 9781 6953 9815 6987
rect 10333 6953 10367 6987
rect 11345 6953 11379 6987
rect 11529 6953 11563 6987
rect 11713 6953 11747 6987
rect 2881 6817 2915 6851
rect 4537 6817 4571 6851
rect 9321 6817 9355 6851
rect 9413 6817 9447 6851
rect 9505 6817 9539 6851
rect 10609 6817 10643 6851
rect 10793 6817 10827 6851
rect 2789 6749 2823 6783
rect 3157 6749 3191 6783
rect 4353 6749 4387 6783
rect 4629 6749 4663 6783
rect 6561 6749 6595 6783
rect 6745 6749 6779 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 8309 6749 8343 6783
rect 9597 6749 9631 6783
rect 10057 6749 10091 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 11437 6749 11471 6783
rect 2697 6681 2731 6715
rect 9781 6681 9815 6715
rect 11681 6681 11715 6715
rect 11897 6681 11931 6715
rect 2329 6613 2363 6647
rect 3341 6613 3375 6647
rect 4721 6613 4755 6647
rect 7665 6613 7699 6647
rect 9965 6613 9999 6647
rect 10977 6613 11011 6647
rect 3893 6409 3927 6443
rect 8493 6409 8527 6443
rect 10609 6409 10643 6443
rect 11253 6409 11287 6443
rect 4169 6341 4203 6375
rect 10333 6341 10367 6375
rect 10517 6341 10551 6375
rect 10977 6341 11011 6375
rect 2053 6273 2087 6307
rect 4261 6273 4295 6307
rect 8677 6273 8711 6307
rect 10149 6273 10183 6307
rect 10793 6273 10827 6307
rect 11069 6273 11103 6307
rect 11161 6273 11195 6307
rect 11345 6273 11379 6307
rect 11713 6273 11747 6307
rect 2145 6205 2179 6239
rect 2421 6205 2455 6239
rect 11897 6137 11931 6171
rect 1869 6069 1903 6103
rect 2881 5865 2915 5899
rect 8769 5865 8803 5899
rect 10701 5865 10735 5899
rect 11805 5865 11839 5899
rect 2789 5797 2823 5831
rect 4261 5797 4295 5831
rect 6377 5797 6411 5831
rect 1409 5729 1443 5763
rect 3433 5729 3467 5763
rect 7297 5729 7331 5763
rect 1676 5661 1710 5695
rect 5549 5661 5583 5695
rect 5917 5661 5951 5695
rect 7021 5661 7055 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 11989 5661 12023 5695
rect 5825 5593 5859 5627
rect 6377 5593 6411 5627
rect 5641 5525 5675 5559
rect 5825 5321 5859 5355
rect 6377 5321 6411 5355
rect 7941 5321 7975 5355
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 6561 5185 6595 5219
rect 7849 5185 7883 5219
rect 11989 5185 12023 5219
rect 3709 5117 3743 5151
rect 3985 5117 4019 5151
rect 5733 5117 5767 5151
rect 6745 5117 6779 5151
rect 11805 4981 11839 5015
rect 4813 4777 4847 4811
rect 9873 4777 9907 4811
rect 10333 4777 10367 4811
rect 4629 4709 4663 4743
rect 8953 4709 8987 4743
rect 9505 4641 9539 4675
rect 10241 4641 10275 4675
rect 4537 4573 4571 4607
rect 4997 4573 5031 4607
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 9137 4573 9171 4607
rect 10057 4573 10091 4607
rect 10517 4573 10551 4607
rect 5089 4505 5123 4539
rect 5181 4505 5215 4539
rect 9229 4505 9263 4539
rect 10333 4505 10367 4539
rect 11253 4505 11287 4539
rect 9321 4437 9355 4471
rect 2789 4233 2823 4267
rect 8493 4233 8527 4267
rect 9597 4233 9631 4267
rect 8125 4165 8159 4199
rect 2697 4097 2731 4131
rect 3893 4097 3927 4131
rect 5549 4097 5583 4131
rect 6929 4097 6963 4131
rect 7113 4097 7147 4131
rect 7297 4097 7331 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 7665 4097 7699 4131
rect 8309 4097 8343 4131
rect 8585 4097 8619 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10609 4097 10643 4131
rect 11161 4097 11195 4131
rect 11529 4097 11563 4131
rect 11621 4097 11655 4131
rect 2881 4029 2915 4063
rect 3617 4029 3651 4063
rect 5825 4029 5859 4063
rect 7941 4029 7975 4063
rect 10425 4029 10459 4063
rect 5641 3961 5675 3995
rect 8309 3961 8343 3995
rect 11069 3961 11103 3995
rect 2329 3893 2363 3927
rect 5733 3893 5767 3927
rect 7389 3893 7423 3927
rect 11529 3893 11563 3927
rect 11897 3893 11931 3927
rect 3617 3689 3651 3723
rect 3985 3689 4019 3723
rect 7113 3689 7147 3723
rect 7757 3689 7791 3723
rect 8953 3689 8987 3723
rect 9597 3689 9631 3723
rect 10149 3689 10183 3723
rect 8677 3621 8711 3655
rect 11713 3621 11747 3655
rect 1869 3553 1903 3587
rect 6469 3553 6503 3587
rect 6561 3553 6595 3587
rect 6653 3553 6687 3587
rect 9965 3553 9999 3587
rect 1777 3485 1811 3519
rect 3893 3485 3927 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 5825 3485 5859 3519
rect 5917 3485 5951 3519
rect 6745 3485 6779 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 7481 3485 7515 3519
rect 7573 3485 7607 3519
rect 7849 3485 7883 3519
rect 7941 3485 7975 3519
rect 8585 3485 8619 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 9505 3485 9539 3519
rect 9781 3485 9815 3519
rect 10057 3485 10091 3519
rect 10241 3485 10275 3519
rect 10701 3485 10735 3519
rect 2145 3417 2179 3451
rect 6193 3417 6227 3451
rect 9321 3417 9355 3451
rect 11897 3417 11931 3451
rect 1593 3349 1627 3383
rect 6285 3349 6319 3383
rect 7297 3349 7331 3383
rect 8033 3349 8067 3383
rect 2881 3145 2915 3179
rect 3709 3145 3743 3179
rect 8769 3145 8803 3179
rect 9873 3145 9907 3179
rect 4445 3077 4479 3111
rect 7297 3077 7331 3111
rect 1409 3009 1443 3043
rect 1676 3009 1710 3043
rect 3801 3009 3835 3043
rect 4169 3009 4203 3043
rect 7021 3009 7055 3043
rect 9781 3009 9815 3043
rect 9965 3009 9999 3043
rect 10701 3009 10735 3043
rect 3433 2941 3467 2975
rect 5917 2941 5951 2975
rect 10609 2941 10643 2975
rect 2789 2873 2823 2907
rect 10333 2873 10367 2907
rect 5181 2601 5215 2635
rect 6101 2601 6135 2635
rect 5089 2397 5123 2431
rect 5917 2397 5951 2431
rect 6837 2397 6871 2431
rect 7481 2397 7515 2431
rect 8125 2397 8159 2431
rect 6653 2261 6687 2295
rect 7297 2261 7331 2295
rect 7941 2261 7975 2295
<< metal1 >>
rect 1104 13082 12328 13104
rect 1104 13030 3013 13082
rect 3065 13030 3077 13082
rect 3129 13030 3141 13082
rect 3193 13030 3205 13082
rect 3257 13030 3269 13082
rect 3321 13030 5819 13082
rect 5871 13030 5883 13082
rect 5935 13030 5947 13082
rect 5999 13030 6011 13082
rect 6063 13030 6075 13082
rect 6127 13030 8625 13082
rect 8677 13030 8689 13082
rect 8741 13030 8753 13082
rect 8805 13030 8817 13082
rect 8869 13030 8881 13082
rect 8933 13030 11431 13082
rect 11483 13030 11495 13082
rect 11547 13030 11559 13082
rect 11611 13030 11623 13082
rect 11675 13030 11687 13082
rect 11739 13030 12328 13082
rect 1104 13008 12328 13030
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5776 12940 5917 12968
rect 5776 12928 5782 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 6512 12872 6561 12900
rect 6512 12860 6518 12872
rect 6549 12869 6561 12872
rect 6595 12869 6607 12903
rect 6549 12863 6607 12869
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5592 12804 5825 12832
rect 5592 12792 5598 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 7156 12804 7205 12832
rect 7156 12792 7162 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 7800 12804 7849 12832
rect 7800 12792 7806 12804
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8444 12804 8677 12832
rect 8444 12792 8450 12804
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 7377 12631 7435 12637
rect 7377 12597 7389 12631
rect 7423 12628 7435 12631
rect 7558 12628 7564 12640
rect 7423 12600 7564 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 8021 12631 8079 12637
rect 8021 12597 8033 12631
rect 8067 12628 8079 12631
rect 8294 12628 8300 12640
rect 8067 12600 8300 12628
rect 8067 12597 8079 12600
rect 8021 12591 8079 12597
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 8478 12588 8484 12640
rect 8536 12588 8542 12640
rect 1104 12538 12328 12560
rect 1104 12486 2353 12538
rect 2405 12486 2417 12538
rect 2469 12486 2481 12538
rect 2533 12486 2545 12538
rect 2597 12486 2609 12538
rect 2661 12486 5159 12538
rect 5211 12486 5223 12538
rect 5275 12486 5287 12538
rect 5339 12486 5351 12538
rect 5403 12486 5415 12538
rect 5467 12486 7965 12538
rect 8017 12486 8029 12538
rect 8081 12486 8093 12538
rect 8145 12486 8157 12538
rect 8209 12486 8221 12538
rect 8273 12486 10771 12538
rect 10823 12486 10835 12538
rect 10887 12486 10899 12538
rect 10951 12486 10963 12538
rect 11015 12486 11027 12538
rect 11079 12486 12328 12538
rect 1104 12464 12328 12486
rect 6178 12316 6184 12368
rect 6236 12356 6242 12368
rect 10321 12359 10379 12365
rect 10321 12356 10333 12359
rect 6236 12328 10333 12356
rect 6236 12316 6242 12328
rect 10321 12325 10333 12328
rect 10367 12325 10379 12359
rect 10321 12319 10379 12325
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 3605 12291 3663 12297
rect 3605 12288 3617 12291
rect 2648 12260 3617 12288
rect 2648 12248 2654 12260
rect 3605 12257 3617 12260
rect 3651 12257 3663 12291
rect 3605 12251 3663 12257
rect 6365 12291 6423 12297
rect 6365 12257 6377 12291
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12288 6699 12291
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 6687 12260 7297 12288
rect 6687 12257 6699 12260
rect 6641 12251 6699 12257
rect 7285 12257 7297 12260
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 4982 12180 4988 12232
rect 5040 12220 5046 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5040 12192 6285 12220
rect 5040 12180 5046 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 1578 12112 1584 12164
rect 1636 12112 1642 12164
rect 2314 12112 2320 12164
rect 2372 12112 2378 12164
rect 3329 12155 3387 12161
rect 3329 12121 3341 12155
rect 3375 12152 3387 12155
rect 4522 12152 4528 12164
rect 3375 12124 4528 12152
rect 3375 12121 3387 12124
rect 3329 12115 3387 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 5353 12155 5411 12161
rect 5353 12121 5365 12155
rect 5399 12152 5411 12155
rect 5534 12152 5540 12164
rect 5399 12124 5540 12152
rect 5399 12121 5411 12124
rect 5353 12115 5411 12121
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 6380 12152 6408 12251
rect 7374 12180 7380 12232
rect 7432 12180 7438 12232
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12220 8079 12223
rect 8294 12220 8300 12232
rect 8067 12192 8300 12220
rect 8067 12189 8079 12192
rect 8021 12183 8079 12189
rect 7558 12152 7564 12164
rect 6380 12124 7564 12152
rect 7558 12112 7564 12124
rect 7616 12112 7622 12164
rect 7852 12152 7880 12183
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 10318 12220 10324 12232
rect 10275 12192 10324 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 10318 12180 10324 12192
rect 10376 12220 10382 12232
rect 10505 12223 10563 12229
rect 10505 12220 10517 12223
rect 10376 12192 10517 12220
rect 10376 12180 10382 12192
rect 10505 12189 10517 12192
rect 10551 12189 10563 12223
rect 10505 12183 10563 12189
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12220 10747 12223
rect 11238 12220 11244 12232
rect 10735 12192 11244 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 8386 12152 8392 12164
rect 7668 12124 8392 12152
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 5626 12084 5632 12096
rect 5307 12056 5632 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 5626 12044 5632 12056
rect 5684 12084 5690 12096
rect 7668 12084 7696 12124
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 9858 12112 9864 12164
rect 9916 12112 9922 12164
rect 10045 12155 10103 12161
rect 10045 12121 10057 12155
rect 10091 12121 10103 12155
rect 10045 12115 10103 12121
rect 5684 12056 7696 12084
rect 5684 12044 5690 12056
rect 7742 12044 7748 12096
rect 7800 12044 7806 12096
rect 7926 12044 7932 12096
rect 7984 12044 7990 12096
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 9306 12084 9312 12096
rect 8168 12056 9312 12084
rect 8168 12044 8174 12056
rect 9306 12044 9312 12056
rect 9364 12084 9370 12096
rect 10060 12084 10088 12115
rect 9364 12056 10088 12084
rect 9364 12044 9370 12056
rect 1104 11994 12328 12016
rect 1104 11942 3013 11994
rect 3065 11942 3077 11994
rect 3129 11942 3141 11994
rect 3193 11942 3205 11994
rect 3257 11942 3269 11994
rect 3321 11942 5819 11994
rect 5871 11942 5883 11994
rect 5935 11942 5947 11994
rect 5999 11942 6011 11994
rect 6063 11942 6075 11994
rect 6127 11942 8625 11994
rect 8677 11942 8689 11994
rect 8741 11942 8753 11994
rect 8805 11942 8817 11994
rect 8869 11942 8881 11994
rect 8933 11942 11431 11994
rect 11483 11942 11495 11994
rect 11547 11942 11559 11994
rect 11611 11942 11623 11994
rect 11675 11942 11687 11994
rect 11739 11942 12328 11994
rect 1104 11920 12328 11942
rect 2314 11840 2320 11892
rect 2372 11880 2378 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2372 11852 2421 11880
rect 2372 11840 2378 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 5534 11880 5540 11892
rect 4387 11852 5540 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 8665 11883 8723 11889
rect 8665 11880 8677 11883
rect 7432 11852 8677 11880
rect 7432 11840 7438 11852
rect 8665 11849 8677 11852
rect 8711 11880 8723 11883
rect 8711 11852 8892 11880
rect 8711 11849 8723 11852
rect 8665 11843 8723 11849
rect 2774 11812 2780 11824
rect 2332 11784 2780 11812
rect 2332 11753 2360 11784
rect 2774 11772 2780 11784
rect 2832 11772 2838 11824
rect 3326 11772 3332 11824
rect 3384 11772 3390 11824
rect 6178 11812 6184 11824
rect 5828 11784 6184 11812
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 2590 11704 2596 11756
rect 2648 11704 2654 11756
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 2869 11679 2927 11685
rect 2869 11645 2881 11679
rect 2915 11676 2927 11679
rect 4525 11679 4583 11685
rect 4525 11676 4537 11679
rect 2915 11648 4537 11676
rect 2915 11645 2927 11648
rect 2869 11639 2927 11645
rect 4525 11645 4537 11648
rect 4571 11645 4583 11679
rect 4724 11676 4752 11707
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 4985 11747 5043 11753
rect 4985 11744 4997 11747
rect 4948 11716 4997 11744
rect 4948 11704 4954 11716
rect 4985 11713 4997 11716
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5534 11744 5540 11756
rect 5215 11716 5540 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 5828 11753 5856 11784
rect 6178 11772 6184 11784
rect 6236 11772 6242 11824
rect 7926 11772 7932 11824
rect 7984 11812 7990 11824
rect 7984 11784 8800 11812
rect 7984 11772 7990 11784
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 6362 11744 6368 11756
rect 5951 11716 6368 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 4724 11648 5457 11676
rect 4525 11639 4583 11645
rect 5445 11645 5457 11648
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 5644 11608 5672 11707
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 7208 11716 7696 11744
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 7208 11676 7236 11716
rect 5767 11648 7236 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 7282 11636 7288 11688
rect 7340 11636 7346 11688
rect 7374 11636 7380 11688
rect 7432 11636 7438 11688
rect 7466 11636 7472 11688
rect 7524 11636 7530 11688
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11645 7619 11679
rect 7668 11676 7696 11716
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 7800 11716 8217 11744
rect 7800 11704 7806 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 8772 11753 8800 11784
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8444 11716 8493 11744
rect 8444 11704 8450 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8864 11744 8892 11852
rect 9306 11840 9312 11892
rect 9364 11840 9370 11892
rect 9858 11840 9864 11892
rect 9916 11840 9922 11892
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8864 11716 8953 11744
rect 8757 11707 8815 11713
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9539 11716 9781 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 7668 11648 7972 11676
rect 7561 11639 7619 11645
rect 6178 11608 6184 11620
rect 5644 11580 6184 11608
rect 6178 11568 6184 11580
rect 6236 11608 6242 11620
rect 6638 11608 6644 11620
rect 6236 11580 6644 11608
rect 6236 11568 6242 11580
rect 6638 11568 6644 11580
rect 6696 11568 6702 11620
rect 7576 11608 7604 11639
rect 7837 11611 7895 11617
rect 7837 11608 7849 11611
rect 7576 11580 7849 11608
rect 7837 11577 7849 11580
rect 7883 11577 7895 11611
rect 7944 11608 7972 11648
rect 8110 11636 8116 11688
rect 8168 11636 8174 11688
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 9508 11676 9536 11707
rect 8895 11648 9536 11676
rect 9677 11679 9735 11685
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 9858 11676 9864 11688
rect 9723 11648 9864 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 9858 11636 9864 11648
rect 9916 11676 9922 11688
rect 9968 11676 9996 11707
rect 10134 11704 10140 11756
rect 10192 11704 10198 11756
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 9916 11648 9996 11676
rect 10612 11676 10640 11707
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 10744 11716 10793 11744
rect 10744 11704 10750 11716
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11146 11744 11152 11756
rect 11103 11716 11152 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11330 11676 11336 11688
rect 10612 11648 11336 11676
rect 9916 11636 9922 11648
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 8386 11608 8392 11620
rect 7944 11580 8392 11608
rect 7837 11571 7895 11577
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 8220 11549 8248 11580
rect 8386 11568 8392 11580
rect 8444 11608 8450 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 8444 11580 10149 11608
rect 8444 11568 8450 11580
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 10137 11571 10195 11577
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 4764 11512 7757 11540
rect 4764 11500 4770 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 8205 11543 8263 11549
rect 8205 11509 8217 11543
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 1104 11450 12328 11472
rect 1104 11398 2353 11450
rect 2405 11398 2417 11450
rect 2469 11398 2481 11450
rect 2533 11398 2545 11450
rect 2597 11398 2609 11450
rect 2661 11398 5159 11450
rect 5211 11398 5223 11450
rect 5275 11398 5287 11450
rect 5339 11398 5351 11450
rect 5403 11398 5415 11450
rect 5467 11398 7965 11450
rect 8017 11398 8029 11450
rect 8081 11398 8093 11450
rect 8145 11398 8157 11450
rect 8209 11398 8221 11450
rect 8273 11398 10771 11450
rect 10823 11398 10835 11450
rect 10887 11398 10899 11450
rect 10951 11398 10963 11450
rect 11015 11398 11027 11450
rect 11079 11398 12328 11450
rect 1104 11376 12328 11398
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 3326 11336 3332 11348
rect 3283 11308 3332 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 4522 11296 4528 11348
rect 4580 11296 4586 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 7006 11336 7012 11348
rect 4948 11308 7012 11336
rect 4948 11296 4954 11308
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 2774 11268 2780 11280
rect 1627 11240 2780 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 2746 11228 2780 11240
rect 2832 11228 2838 11280
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 2746 11132 2774 11228
rect 4982 11160 4988 11212
rect 5040 11160 5046 11212
rect 5276 11209 5304 11308
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7524 11308 7665 11336
rect 7524 11296 7530 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7653 11299 7711 11305
rect 7745 11339 7803 11345
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 8386 11336 8392 11348
rect 7791 11308 8392 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 11238 11296 11244 11348
rect 11296 11296 11302 11348
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 5460 11240 10057 11268
rect 5261 11203 5319 11209
rect 5460 11208 5488 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 11388 11240 11652 11268
rect 11388 11228 11394 11240
rect 5261 11169 5273 11203
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5368 11180 5488 11208
rect 7561 11203 7619 11209
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 2746 11104 3157 11132
rect 3145 11101 3157 11104
rect 3191 11132 3203 11135
rect 3418 11132 3424 11144
rect 3191 11104 3424 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 4706 11092 4712 11144
rect 4764 11092 4770 11144
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5368 11132 5396 11180
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7650 11200 7656 11212
rect 7607 11172 7656 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 11624 11209 11652 11240
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 7760 11172 10333 11200
rect 5215 11104 5396 11132
rect 5445 11135 5503 11141
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5445 11101 5457 11135
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 4982 11064 4988 11076
rect 1636 11036 4988 11064
rect 1636 11024 1642 11036
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 5460 11064 5488 11095
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 6546 11132 6552 11144
rect 5951 11104 6552 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 7760 11132 7788 11172
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 10321 11163 10379 11169
rect 10428 11172 10517 11200
rect 6696 11104 7788 11132
rect 6696 11092 6702 11104
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 10428 11141 10456 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 10505 11163 10563 11169
rect 10980 11172 11529 11200
rect 10980 11144 11008 11172
rect 11517 11169 11529 11172
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11169 11667 11203
rect 11609 11163 11667 11169
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 11204 11104 11437 11132
rect 11204 11092 11210 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 5813 11067 5871 11073
rect 5813 11064 5825 11067
rect 5460 11036 5825 11064
rect 5813 11033 5825 11036
rect 5859 11033 5871 11067
rect 5813 11027 5871 11033
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 8386 11064 8392 11076
rect 7432 11036 8392 11064
rect 7432 11024 7438 11036
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 10888 11064 10916 11092
rect 11716 11064 11744 11095
rect 10888 11036 11744 11064
rect 5350 10956 5356 11008
rect 5408 10956 5414 11008
rect 1104 10906 12328 10928
rect 1104 10854 3013 10906
rect 3065 10854 3077 10906
rect 3129 10854 3141 10906
rect 3193 10854 3205 10906
rect 3257 10854 3269 10906
rect 3321 10854 5819 10906
rect 5871 10854 5883 10906
rect 5935 10854 5947 10906
rect 5999 10854 6011 10906
rect 6063 10854 6075 10906
rect 6127 10854 8625 10906
rect 8677 10854 8689 10906
rect 8741 10854 8753 10906
rect 8805 10854 8817 10906
rect 8869 10854 8881 10906
rect 8933 10854 11431 10906
rect 11483 10854 11495 10906
rect 11547 10854 11559 10906
rect 11611 10854 11623 10906
rect 11675 10854 11687 10906
rect 11739 10854 12328 10906
rect 1104 10832 12328 10854
rect 5350 10792 5356 10804
rect 1688 10764 5356 10792
rect 1688 10733 1716 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6362 10752 6368 10804
rect 6420 10752 6426 10804
rect 8128 10764 8708 10792
rect 1673 10727 1731 10733
rect 1673 10693 1685 10727
rect 1719 10693 1731 10727
rect 3329 10727 3387 10733
rect 3329 10724 3341 10727
rect 2898 10696 3341 10724
rect 1673 10687 1731 10693
rect 3329 10693 3341 10696
rect 3375 10693 3387 10727
rect 6914 10724 6920 10736
rect 3329 10687 3387 10693
rect 5368 10696 6920 10724
rect 3418 10616 3424 10668
rect 3476 10616 3482 10668
rect 5368 10665 5396 10696
rect 6914 10684 6920 10696
rect 6972 10724 6978 10736
rect 8128 10724 8156 10764
rect 8478 10724 8484 10736
rect 6972 10696 8156 10724
rect 8220 10696 8484 10724
rect 6972 10684 6978 10696
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5000 10628 5365 10656
rect 1394 10548 1400 10600
rect 1452 10548 1458 10600
rect 3145 10591 3203 10597
rect 3145 10557 3157 10591
rect 3191 10588 3203 10591
rect 5000 10588 5028 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 8220 10665 8248 10696
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 8680 10733 8708 10764
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 10962 10792 10968 10804
rect 10744 10764 10968 10792
rect 10744 10752 10750 10764
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 8665 10727 8723 10733
rect 8665 10693 8677 10727
rect 8711 10693 8723 10727
rect 8665 10687 8723 10693
rect 10410 10684 10416 10736
rect 10468 10724 10474 10736
rect 10597 10727 10655 10733
rect 10597 10724 10609 10727
rect 10468 10696 10609 10724
rect 10468 10684 10474 10696
rect 10597 10693 10609 10696
rect 10643 10693 10655 10727
rect 11241 10727 11299 10733
rect 11241 10724 11253 10727
rect 10597 10687 10655 10693
rect 10796 10696 11253 10724
rect 10796 10668 10824 10696
rect 11241 10693 11253 10696
rect 11287 10693 11299 10727
rect 11241 10687 11299 10693
rect 8113 10659 8171 10665
rect 8113 10656 8125 10659
rect 7616 10628 8125 10656
rect 7616 10616 7622 10628
rect 8113 10625 8125 10628
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 8570 10656 8576 10668
rect 8435 10628 8576 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 9858 10656 9864 10668
rect 8895 10628 9864 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 11057 10659 11115 10665
rect 11057 10625 11069 10659
rect 11103 10656 11115 10659
rect 11146 10656 11152 10668
rect 11103 10628 11152 10656
rect 11103 10625 11115 10628
rect 11057 10619 11115 10625
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11330 10616 11336 10668
rect 11388 10616 11394 10668
rect 3191 10560 5028 10588
rect 5077 10591 5135 10597
rect 3191 10557 3203 10560
rect 3145 10551 3203 10557
rect 5077 10557 5089 10591
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 5092 10520 5120 10551
rect 5534 10548 5540 10600
rect 5592 10548 5598 10600
rect 6822 10548 6828 10600
rect 6880 10548 6886 10600
rect 10134 10548 10140 10600
rect 10192 10588 10198 10600
rect 10689 10591 10747 10597
rect 10689 10588 10701 10591
rect 10192 10560 10701 10588
rect 10192 10548 10198 10560
rect 10689 10557 10701 10560
rect 10735 10588 10747 10591
rect 10870 10588 10876 10600
rect 10735 10560 10876 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 5718 10520 5724 10532
rect 5092 10492 5724 10520
rect 5718 10480 5724 10492
rect 5776 10520 5782 10532
rect 5902 10520 5908 10532
rect 5776 10492 5908 10520
rect 5776 10480 5782 10492
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 5997 10523 6055 10529
rect 5997 10489 6009 10523
rect 6043 10520 6055 10523
rect 6733 10523 6791 10529
rect 6733 10520 6745 10523
rect 6043 10492 6745 10520
rect 6043 10489 6055 10492
rect 5997 10483 6055 10489
rect 6733 10489 6745 10492
rect 6779 10489 6791 10523
rect 6733 10483 6791 10489
rect 7929 10523 7987 10529
rect 7929 10489 7941 10523
rect 7975 10520 7987 10523
rect 9582 10520 9588 10532
rect 7975 10492 9588 10520
rect 7975 10489 7987 10492
rect 7929 10483 7987 10489
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 8294 10412 8300 10464
rect 8352 10412 8358 10464
rect 1104 10362 12328 10384
rect 1104 10310 2353 10362
rect 2405 10310 2417 10362
rect 2469 10310 2481 10362
rect 2533 10310 2545 10362
rect 2597 10310 2609 10362
rect 2661 10310 5159 10362
rect 5211 10310 5223 10362
rect 5275 10310 5287 10362
rect 5339 10310 5351 10362
rect 5403 10310 5415 10362
rect 5467 10310 7965 10362
rect 8017 10310 8029 10362
rect 8081 10310 8093 10362
rect 8145 10310 8157 10362
rect 8209 10310 8221 10362
rect 8273 10310 10771 10362
rect 10823 10310 10835 10362
rect 10887 10310 10899 10362
rect 10951 10310 10963 10362
rect 11015 10310 11027 10362
rect 11079 10310 12328 10362
rect 1104 10288 12328 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 1489 10251 1547 10257
rect 1489 10248 1501 10251
rect 1360 10220 1501 10248
rect 1360 10208 1366 10220
rect 1489 10217 1501 10220
rect 1535 10217 1547 10251
rect 1489 10211 1547 10217
rect 4985 10251 5043 10257
rect 4985 10217 4997 10251
rect 5031 10248 5043 10251
rect 5074 10248 5080 10260
rect 5031 10220 5080 10248
rect 5031 10217 5043 10220
rect 4985 10211 5043 10217
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 10134 10208 10140 10260
rect 10192 10208 10198 10260
rect 5552 10180 5580 10208
rect 5368 10152 5580 10180
rect 1578 10004 1584 10056
rect 1636 10044 1642 10056
rect 5368 10053 5396 10152
rect 5994 10140 6000 10192
rect 6052 10180 6058 10192
rect 6052 10152 8248 10180
rect 6052 10140 6058 10152
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 5460 10084 6101 10112
rect 5460 10053 5488 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 6089 10075 6147 10081
rect 1673 10047 1731 10053
rect 1673 10044 1685 10047
rect 1636 10016 1685 10044
rect 1636 10004 1642 10016
rect 1673 10013 1685 10016
rect 1719 10013 1731 10047
rect 5169 10047 5227 10053
rect 5169 10044 5181 10047
rect 1673 10007 1731 10013
rect 5000 10016 5181 10044
rect 5000 9908 5028 10016
rect 5169 10013 5181 10016
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5994 10044 6000 10056
rect 5767 10016 6000 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5074 9936 5080 9988
rect 5132 9976 5138 9988
rect 5736 9976 5764 10007
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 8220 10053 8248 10152
rect 9122 10140 9128 10192
rect 9180 10180 9186 10192
rect 9401 10183 9459 10189
rect 9401 10180 9413 10183
rect 9180 10152 9413 10180
rect 9180 10140 9186 10152
rect 9401 10149 9413 10152
rect 9447 10149 9459 10183
rect 9401 10143 9459 10149
rect 11793 10183 11851 10189
rect 11793 10149 11805 10183
rect 11839 10149 11851 10183
rect 11793 10143 11851 10149
rect 9858 10072 9864 10124
rect 9916 10072 9922 10124
rect 6181 10047 6239 10053
rect 6181 10046 6193 10047
rect 6104 10018 6193 10046
rect 5132 9948 5764 9976
rect 5905 9979 5963 9985
rect 5132 9936 5138 9948
rect 5905 9945 5917 9979
rect 5951 9976 5963 9979
rect 6104 9976 6132 10018
rect 6181 10013 6193 10018
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 8205 10007 8263 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8478 10044 8484 10056
rect 8435 10016 8484 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 11808 10044 11836 10143
rect 9416 10016 11836 10044
rect 9416 9988 9444 10016
rect 11974 10004 11980 10056
rect 12032 10004 12038 10056
rect 6362 9976 6368 9988
rect 5951 9948 6368 9976
rect 5951 9945 5963 9948
rect 5905 9939 5963 9945
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 8570 9936 8576 9988
rect 8628 9976 8634 9988
rect 9398 9976 9404 9988
rect 8628 9948 9404 9976
rect 8628 9936 8634 9948
rect 9398 9936 9404 9948
rect 9456 9936 9462 9988
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 9508 9948 9965 9976
rect 6454 9908 6460 9920
rect 5000 9880 6460 9908
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 9306 9908 9312 9920
rect 8343 9880 9312 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 9306 9868 9312 9880
rect 9364 9908 9370 9920
rect 9508 9908 9536 9948
rect 9953 9945 9965 9948
rect 9999 9945 10011 9979
rect 9953 9939 10011 9945
rect 9364 9880 9536 9908
rect 9364 9868 9370 9880
rect 1104 9818 12328 9840
rect 1104 9766 3013 9818
rect 3065 9766 3077 9818
rect 3129 9766 3141 9818
rect 3193 9766 3205 9818
rect 3257 9766 3269 9818
rect 3321 9766 5819 9818
rect 5871 9766 5883 9818
rect 5935 9766 5947 9818
rect 5999 9766 6011 9818
rect 6063 9766 6075 9818
rect 6127 9766 8625 9818
rect 8677 9766 8689 9818
rect 8741 9766 8753 9818
rect 8805 9766 8817 9818
rect 8869 9766 8881 9818
rect 8933 9766 11431 9818
rect 11483 9766 11495 9818
rect 11547 9766 11559 9818
rect 11611 9766 11623 9818
rect 11675 9766 11687 9818
rect 11739 9766 12328 9818
rect 1104 9744 12328 9766
rect 9858 9704 9864 9716
rect 9232 9676 9864 9704
rect 7282 9596 7288 9648
rect 7340 9596 7346 9648
rect 9232 9645 9260 9676
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 9217 9639 9275 9645
rect 9217 9605 9229 9639
rect 9263 9605 9275 9639
rect 9217 9599 9275 9605
rect 9306 9596 9312 9648
rect 9364 9596 9370 9648
rect 2774 9528 2780 9580
rect 2832 9528 2838 9580
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 6822 9568 6828 9580
rect 6512 9540 6828 9568
rect 6512 9528 6518 9540
rect 6822 9528 6828 9540
rect 6880 9568 6886 9580
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6880 9540 7021 9568
rect 6880 9528 6886 9540
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 9398 9528 9404 9580
rect 9456 9568 9462 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9456 9540 9597 9568
rect 9456 9528 9462 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 1394 9460 1400 9512
rect 1452 9460 1458 9512
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 2740 9472 3249 9500
rect 2740 9460 2746 9472
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 3237 9463 3295 9469
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 6604 9472 7297 9500
rect 6604 9460 6610 9472
rect 7285 9469 7297 9472
rect 7331 9500 7343 9503
rect 7466 9500 7472 9512
rect 7331 9472 7472 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 9180 9472 9689 9500
rect 9180 9460 9186 9472
rect 9677 9469 9689 9472
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 1412 9364 1440 9460
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9432 9919 9435
rect 11330 9432 11336 9444
rect 9907 9404 11336 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 11330 9392 11336 9404
rect 11388 9392 11394 9444
rect 2682 9364 2688 9376
rect 1412 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 5534 9364 5540 9376
rect 3191 9336 5540 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 7101 9367 7159 9373
rect 7101 9364 7113 9367
rect 5960 9336 7113 9364
rect 5960 9324 5966 9336
rect 7101 9333 7113 9336
rect 7147 9333 7159 9367
rect 7101 9327 7159 9333
rect 1104 9274 12328 9296
rect 1104 9222 2353 9274
rect 2405 9222 2417 9274
rect 2469 9222 2481 9274
rect 2533 9222 2545 9274
rect 2597 9222 2609 9274
rect 2661 9222 5159 9274
rect 5211 9222 5223 9274
rect 5275 9222 5287 9274
rect 5339 9222 5351 9274
rect 5403 9222 5415 9274
rect 5467 9222 7965 9274
rect 8017 9222 8029 9274
rect 8081 9222 8093 9274
rect 8145 9222 8157 9274
rect 8209 9222 8221 9274
rect 8273 9222 10771 9274
rect 10823 9222 10835 9274
rect 10887 9222 10899 9274
rect 10951 9222 10963 9274
rect 11015 9222 11027 9274
rect 11079 9222 12328 9274
rect 1104 9200 12328 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 2409 9163 2467 9169
rect 2409 9160 2421 9163
rect 1728 9132 2421 9160
rect 1728 9120 1734 9132
rect 2409 9129 2421 9132
rect 2455 9129 2467 9163
rect 2409 9123 2467 9129
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2832 9132 2881 9160
rect 2832 9120 2838 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 2869 9123 2927 9129
rect 5902 9120 5908 9172
rect 5960 9120 5966 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 9122 9160 9128 9172
rect 8352 9132 9128 9160
rect 8352 9120 8358 9132
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 10560 9132 11897 9160
rect 10560 9120 10566 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 7745 9095 7803 9101
rect 7745 9092 7757 9095
rect 2608 9064 7757 9092
rect 2608 8965 2636 9064
rect 7745 9061 7757 9064
rect 7791 9061 7803 9095
rect 7745 9055 7803 9061
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 11149 9095 11207 9101
rect 11149 9092 11161 9095
rect 10744 9064 11161 9092
rect 10744 9052 10750 9064
rect 11149 9061 11161 9064
rect 11195 9092 11207 9095
rect 11195 9064 11836 9092
rect 11195 9061 11207 9064
rect 11149 9055 11207 9061
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 3237 9027 3295 9033
rect 3237 9024 3249 9027
rect 2740 8996 3249 9024
rect 2740 8984 2746 8996
rect 3237 8993 3249 8996
rect 3283 8993 3295 9027
rect 3237 8987 3295 8993
rect 5718 8984 5724 9036
rect 5776 8984 5782 9036
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 8297 9027 8355 9033
rect 8297 9024 8309 9027
rect 7524 8996 8309 9024
rect 7524 8984 7530 8996
rect 8297 8993 8309 8996
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 9398 8984 9404 9036
rect 9456 9024 9462 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9456 8996 10057 9024
rect 9456 8984 9462 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2593 8919 2651 8925
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3418 8956 3424 8968
rect 3007 8928 3424 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3418 8916 3424 8928
rect 3476 8956 3482 8968
rect 3786 8956 3792 8968
rect 3476 8928 3792 8956
rect 3476 8916 3482 8928
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 5258 8956 5264 8968
rect 4948 8928 5264 8956
rect 4948 8916 4954 8928
rect 5258 8916 5264 8928
rect 5316 8956 5322 8968
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 5316 8928 5641 8956
rect 5316 8916 5322 8928
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 5629 8919 5687 8925
rect 7392 8928 8953 8956
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 7392 8888 7420 8928
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 10134 8956 10140 8968
rect 8987 8928 10140 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 5592 8860 7420 8888
rect 5592 8848 5598 8860
rect 7466 8848 7472 8900
rect 7524 8848 7530 8900
rect 8113 8891 8171 8897
rect 8113 8857 8125 8891
rect 8159 8888 8171 8891
rect 8294 8888 8300 8900
rect 8159 8860 8300 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7558 8820 7564 8832
rect 7064 8792 7564 8820
rect 7064 8780 7070 8792
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 8202 8780 8208 8832
rect 8260 8780 8266 8832
rect 10505 8823 10563 8829
rect 10505 8789 10517 8823
rect 10551 8820 10563 8823
rect 10980 8820 11008 8919
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11808 8965 11836 9064
rect 11793 8959 11851 8965
rect 11204 8928 11376 8956
rect 11204 8916 11210 8928
rect 11348 8897 11376 8928
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 11333 8891 11391 8897
rect 11333 8857 11345 8891
rect 11379 8857 11391 8891
rect 11333 8851 11391 8857
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8857 11575 8891
rect 11517 8851 11575 8857
rect 11701 8891 11759 8897
rect 11701 8857 11713 8891
rect 11747 8888 11759 8891
rect 11992 8888 12020 8919
rect 11747 8860 12020 8888
rect 11747 8857 11759 8860
rect 11701 8851 11759 8857
rect 11532 8820 11560 8851
rect 10551 8792 11560 8820
rect 10551 8789 10563 8792
rect 10505 8783 10563 8789
rect 1104 8730 12328 8752
rect 1104 8678 3013 8730
rect 3065 8678 3077 8730
rect 3129 8678 3141 8730
rect 3193 8678 3205 8730
rect 3257 8678 3269 8730
rect 3321 8678 5819 8730
rect 5871 8678 5883 8730
rect 5935 8678 5947 8730
rect 5999 8678 6011 8730
rect 6063 8678 6075 8730
rect 6127 8678 8625 8730
rect 8677 8678 8689 8730
rect 8741 8678 8753 8730
rect 8805 8678 8817 8730
rect 8869 8678 8881 8730
rect 8933 8678 11431 8730
rect 11483 8678 11495 8730
rect 11547 8678 11559 8730
rect 11611 8678 11623 8730
rect 11675 8678 11687 8730
rect 11739 8678 12328 8730
rect 1104 8656 12328 8678
rect 2682 8576 2688 8628
rect 2740 8576 2746 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5776 8588 6009 8616
rect 5776 8576 5782 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 6917 8619 6975 8625
rect 6917 8616 6929 8619
rect 6420 8588 6929 8616
rect 6420 8576 6426 8588
rect 6917 8585 6929 8588
rect 6963 8585 6975 8619
rect 6917 8579 6975 8585
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8260 8588 9229 8616
rect 8260 8576 8266 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9217 8579 9275 8585
rect 11882 8576 11888 8628
rect 11940 8576 11946 8628
rect 2700 8548 2728 8576
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 2700 8520 3372 8548
rect 3344 8489 3372 8520
rect 5000 8520 5365 8548
rect 5000 8489 5028 8520
rect 5353 8517 5365 8520
rect 5399 8548 5411 8551
rect 6638 8548 6644 8560
rect 5399 8520 6644 8548
rect 5399 8517 5411 8520
rect 5353 8511 5411 8517
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 9030 8548 9036 8560
rect 8864 8520 9036 8548
rect 3329 8483 3387 8489
rect 1964 8412 1992 8466
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 2958 8412 2964 8424
rect 1964 8384 2964 8412
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3050 8372 3056 8424
rect 3108 8372 3114 8424
rect 1578 8236 1584 8288
rect 1636 8236 1642 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4617 8279 4675 8285
rect 4617 8276 4629 8279
rect 4212 8248 4629 8276
rect 4212 8236 4218 8248
rect 4617 8245 4629 8248
rect 4663 8245 4675 8279
rect 4816 8276 4844 8443
rect 5092 8412 5120 8443
rect 5258 8440 5264 8492
rect 5316 8440 5322 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5828 8452 5917 8480
rect 5644 8412 5672 8440
rect 5092 8384 5672 8412
rect 4893 8347 4951 8353
rect 4893 8313 4905 8347
rect 4939 8344 4951 8347
rect 4939 8316 5488 8344
rect 4939 8313 4951 8316
rect 4893 8307 4951 8313
rect 5074 8276 5080 8288
rect 4816 8248 5080 8276
rect 4617 8239 4675 8245
rect 5074 8236 5080 8248
rect 5132 8276 5138 8288
rect 5353 8279 5411 8285
rect 5353 8276 5365 8279
rect 5132 8248 5365 8276
rect 5132 8236 5138 8248
rect 5353 8245 5365 8248
rect 5399 8245 5411 8279
rect 5460 8276 5488 8316
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 5828 8353 5856 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8480 6147 8483
rect 6730 8480 6736 8492
rect 6135 8452 6736 8480
rect 6135 8449 6147 8452
rect 6089 8443 6147 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 6822 8440 6828 8492
rect 6880 8440 6886 8492
rect 7098 8440 7104 8492
rect 7156 8440 7162 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8864 8489 8892 8520
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 11054 8548 11060 8560
rect 10060 8520 11060 8548
rect 10060 8492 10088 8520
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8444 8452 8861 8480
rect 8444 8440 8450 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8480 8999 8483
rect 10042 8480 10048 8492
rect 8987 8452 10048 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 10192 8452 11713 8480
rect 10192 8440 10198 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6472 8384 6653 8412
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5592 8316 5825 8344
rect 5592 8304 5598 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5813 8307 5871 8313
rect 6472 8276 6500 8384
rect 6641 8381 6653 8384
rect 6687 8412 6699 8415
rect 8294 8412 8300 8424
rect 6687 8384 8300 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 10410 8412 10416 8424
rect 9079 8384 10416 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 8772 8344 8800 8375
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 7147 8316 8800 8344
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 6546 8276 6552 8288
rect 5460 8248 6552 8276
rect 5353 8239 5411 8245
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6638 8236 6644 8288
rect 6696 8236 6702 8288
rect 1104 8186 12328 8208
rect 1104 8134 2353 8186
rect 2405 8134 2417 8186
rect 2469 8134 2481 8186
rect 2533 8134 2545 8186
rect 2597 8134 2609 8186
rect 2661 8134 5159 8186
rect 5211 8134 5223 8186
rect 5275 8134 5287 8186
rect 5339 8134 5351 8186
rect 5403 8134 5415 8186
rect 5467 8134 7965 8186
rect 8017 8134 8029 8186
rect 8081 8134 8093 8186
rect 8145 8134 8157 8186
rect 8209 8134 8221 8186
rect 8273 8134 10771 8186
rect 10823 8134 10835 8186
rect 10887 8134 10899 8186
rect 10951 8134 10963 8186
rect 11015 8134 11027 8186
rect 11079 8134 12328 8186
rect 1104 8112 12328 8134
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 1489 8075 1547 8081
rect 1489 8072 1501 8075
rect 1360 8044 1501 8072
rect 1360 8032 1366 8044
rect 1489 8041 1501 8044
rect 1535 8041 1547 8075
rect 1489 8035 1547 8041
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 3108 8044 3157 8072
rect 3108 8032 3114 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3145 8035 3203 8041
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5442 8072 5448 8084
rect 5040 8044 5448 8072
rect 5040 8032 5046 8044
rect 5442 8032 5448 8044
rect 5500 8072 5506 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5500 8044 5549 8072
rect 5500 8032 5506 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 6822 8032 6828 8084
rect 6880 8032 6886 8084
rect 10410 8032 10416 8084
rect 10468 8032 10474 8084
rect 2958 7964 2964 8016
rect 3016 8004 3022 8016
rect 3881 8007 3939 8013
rect 3881 8004 3893 8007
rect 3016 7976 3893 8004
rect 3016 7964 3022 7976
rect 3881 7973 3893 7976
rect 3927 8004 3939 8007
rect 4062 8004 4068 8016
rect 3927 7976 4068 8004
rect 3927 7973 3939 7976
rect 3881 7967 3939 7973
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 7466 7964 7472 8016
rect 7524 8004 7530 8016
rect 8202 8004 8208 8016
rect 7524 7976 8208 8004
rect 7524 7964 7530 7976
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 4522 7936 4528 7948
rect 3620 7908 4528 7936
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 3620 7877 3648 7908
rect 4522 7896 4528 7908
rect 4580 7936 4586 7948
rect 6178 7936 6184 7948
rect 4580 7908 6184 7936
rect 4580 7896 4586 7908
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 1673 7871 1731 7877
rect 1673 7868 1685 7871
rect 1636 7840 1685 7868
rect 1636 7828 1642 7840
rect 1673 7837 1685 7840
rect 1719 7868 1731 7871
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 1719 7840 2421 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3099 7840 3341 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 4246 7828 4252 7880
rect 4304 7828 4310 7880
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6604 7840 6745 7868
rect 6604 7828 6610 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 10318 7828 10324 7880
rect 10376 7828 10382 7880
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 6457 7803 6515 7809
rect 6457 7769 6469 7803
rect 6503 7800 6515 7803
rect 7098 7800 7104 7812
rect 6503 7772 7104 7800
rect 6503 7769 6515 7772
rect 6457 7763 6515 7769
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 8389 7803 8447 7809
rect 8389 7769 8401 7803
rect 8435 7800 8447 7803
rect 9122 7800 9128 7812
rect 8435 7772 9128 7800
rect 8435 7769 8447 7772
rect 8389 7763 8447 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 3513 7735 3571 7741
rect 3513 7732 3525 7735
rect 2832 7704 3525 7732
rect 2832 7692 2838 7704
rect 3513 7701 3525 7704
rect 3559 7701 3571 7735
rect 3513 7695 3571 7701
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 6822 7732 6828 7744
rect 6604 7704 6828 7732
rect 6604 7692 6610 7704
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 1104 7642 12328 7664
rect 1104 7590 3013 7642
rect 3065 7590 3077 7642
rect 3129 7590 3141 7642
rect 3193 7590 3205 7642
rect 3257 7590 3269 7642
rect 3321 7590 5819 7642
rect 5871 7590 5883 7642
rect 5935 7590 5947 7642
rect 5999 7590 6011 7642
rect 6063 7590 6075 7642
rect 6127 7590 8625 7642
rect 8677 7590 8689 7642
rect 8741 7590 8753 7642
rect 8805 7590 8817 7642
rect 8869 7590 8881 7642
rect 8933 7590 11431 7642
rect 11483 7590 11495 7642
rect 11547 7590 11559 7642
rect 11611 7590 11623 7642
rect 11675 7590 11687 7642
rect 11739 7590 12328 7642
rect 1104 7568 12328 7590
rect 6641 7531 6699 7537
rect 3896 7500 5764 7528
rect 3896 7404 3924 7500
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 4120 7432 4384 7460
rect 4120 7420 4126 7432
rect 3878 7352 3884 7404
rect 3936 7352 3942 7404
rect 4356 7401 4384 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4062 7284 4068 7336
rect 4120 7284 4126 7336
rect 3970 7216 3976 7268
rect 4028 7216 4034 7268
rect 2682 7148 2688 7200
rect 2740 7188 2746 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 2740 7160 3709 7188
rect 2740 7148 2746 7160
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 4172 7188 4200 7355
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4948 7364 5089 7392
rect 4948 7352 4954 7364
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5534 7392 5540 7404
rect 5491 7364 5540 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 5736 7401 5764 7500
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6914 7528 6920 7540
rect 6687 7500 6920 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6914 7488 6920 7500
rect 6972 7528 6978 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 6972 7500 7481 7528
rect 6972 7488 6978 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 7469 7491 7527 7497
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8260 7500 8616 7528
rect 8260 7488 8266 7500
rect 7009 7463 7067 7469
rect 7009 7429 7021 7463
rect 7055 7460 7067 7463
rect 7055 7432 8524 7460
rect 7055 7429 7067 7432
rect 7009 7423 7067 7429
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 6822 7352 6828 7404
rect 6880 7352 6886 7404
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 8202 7392 8208 7404
rect 7331 7364 8208 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 7116 7324 7144 7355
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 6788 7296 7144 7324
rect 8312 7324 8340 7355
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 8496 7401 8524 7432
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7361 8539 7395
rect 8588 7392 8616 7500
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 8720 7500 8984 7528
rect 8720 7488 8726 7500
rect 8956 7469 8984 7500
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10100 7500 10333 7528
rect 10100 7488 10106 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 10502 7488 10508 7540
rect 10560 7488 10566 7540
rect 8941 7463 8999 7469
rect 8941 7429 8953 7463
rect 8987 7429 8999 7463
rect 8941 7423 8999 7429
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8588 7364 8677 7392
rect 8481 7355 8539 7361
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8754 7352 8760 7404
rect 8812 7352 8818 7404
rect 9140 7392 9168 7488
rect 10520 7460 10548 7488
rect 10520 7432 11008 7460
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9140 7364 9413 7392
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9582 7352 9588 7404
rect 9640 7352 9646 7404
rect 10502 7352 10508 7404
rect 10560 7352 10566 7404
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 9766 7324 9772 7336
rect 8312 7296 9772 7324
rect 6788 7284 6794 7296
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10612 7324 10640 7355
rect 10686 7352 10692 7404
rect 10744 7352 10750 7404
rect 10778 7352 10784 7404
rect 10836 7352 10842 7404
rect 10980 7401 11008 7432
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 10468 7296 10640 7324
rect 10468 7284 10474 7296
rect 9217 7259 9275 7265
rect 9217 7256 9229 7259
rect 5644 7228 9229 7256
rect 5644 7188 5672 7228
rect 9217 7225 9229 7228
rect 9263 7225 9275 7259
rect 9217 7219 9275 7225
rect 4172 7160 5672 7188
rect 6181 7191 6239 7197
rect 3697 7151 3755 7157
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 7098 7188 7104 7200
rect 6227 7160 7104 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7892 7160 8033 7188
rect 7892 7148 7898 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 9582 7148 9588 7200
rect 9640 7148 9646 7200
rect 1104 7098 12328 7120
rect 1104 7046 2353 7098
rect 2405 7046 2417 7098
rect 2469 7046 2481 7098
rect 2533 7046 2545 7098
rect 2597 7046 2609 7098
rect 2661 7046 5159 7098
rect 5211 7046 5223 7098
rect 5275 7046 5287 7098
rect 5339 7046 5351 7098
rect 5403 7046 5415 7098
rect 5467 7046 7965 7098
rect 8017 7046 8029 7098
rect 8081 7046 8093 7098
rect 8145 7046 8157 7098
rect 8209 7046 8221 7098
rect 8273 7046 10771 7098
rect 10823 7046 10835 7098
rect 10887 7046 10899 7098
rect 10951 7046 10963 7098
rect 11015 7046 11027 7098
rect 11079 7046 12328 7098
rect 1104 7024 12328 7046
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 6641 6987 6699 6993
rect 6641 6984 6653 6987
rect 6604 6956 6653 6984
rect 6604 6944 6610 6956
rect 6641 6953 6653 6956
rect 6687 6953 6699 6987
rect 6641 6947 6699 6953
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 9125 6987 9183 6993
rect 9125 6984 9137 6987
rect 8444 6956 9137 6984
rect 8444 6944 8450 6956
rect 9125 6953 9137 6956
rect 9171 6953 9183 6987
rect 9674 6984 9680 6996
rect 9125 6947 9183 6953
rect 9324 6956 9680 6984
rect 6178 6916 6184 6928
rect 4632 6888 6184 6916
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2740 6820 2881 6848
rect 2740 6808 2746 6820
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 4522 6808 4528 6860
rect 4580 6808 4586 6860
rect 2774 6740 2780 6792
rect 2832 6740 2838 6792
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3786 6780 3792 6792
rect 3191 6752 3792 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4632 6789 4660 6888
rect 6178 6876 6184 6888
rect 6236 6916 6242 6928
rect 8754 6916 8760 6928
rect 6236 6888 8760 6916
rect 6236 6876 6242 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 6638 6848 6644 6860
rect 6564 6820 6644 6848
rect 6564 6789 6592 6820
rect 6638 6808 6644 6820
rect 6696 6848 6702 6860
rect 9324 6857 9352 6956
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 9766 6944 9772 6996
rect 9824 6944 9830 6996
rect 10318 6944 10324 6996
rect 10376 6944 10382 6996
rect 10686 6944 10692 6996
rect 10744 6984 10750 6996
rect 11333 6987 11391 6993
rect 11333 6984 11345 6987
rect 10744 6956 11345 6984
rect 10744 6944 10750 6956
rect 9950 6916 9956 6928
rect 9416 6888 9956 6916
rect 9416 6857 9444 6888
rect 9950 6876 9956 6888
rect 10008 6916 10014 6928
rect 10410 6916 10416 6928
rect 10008 6888 10416 6916
rect 10008 6876 10014 6888
rect 10410 6876 10416 6888
rect 10468 6916 10474 6928
rect 10468 6888 10640 6916
rect 10468 6876 10474 6888
rect 9309 6851 9367 6857
rect 6696 6820 8340 6848
rect 6696 6808 6702 6820
rect 8312 6792 8340 6820
rect 9309 6817 9321 6851
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9766 6848 9772 6860
rect 9539 6820 9772 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 10612 6857 10640 6888
rect 10796 6857 10824 6956
rect 11333 6953 11345 6956
rect 11379 6984 11391 6987
rect 11517 6987 11575 6993
rect 11517 6984 11529 6987
rect 11379 6956 11529 6984
rect 11379 6953 11391 6956
rect 11333 6947 11391 6953
rect 11517 6953 11529 6956
rect 11563 6953 11575 6987
rect 11517 6947 11575 6953
rect 11701 6987 11759 6993
rect 11701 6953 11713 6987
rect 11747 6953 11759 6987
rect 11701 6947 11759 6953
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 11716 6916 11744 6947
rect 10928 6888 11744 6916
rect 10928 6876 10934 6888
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4028 6752 4353 6780
rect 4028 6740 4034 6752
rect 4341 6749 4353 6752
rect 4387 6780 4399 6783
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4387 6752 4629 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 7834 6740 7840 6792
rect 7892 6740 7898 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 2685 6715 2743 6721
rect 2685 6681 2697 6715
rect 2731 6712 2743 6715
rect 2866 6712 2872 6724
rect 2731 6684 2872 6712
rect 2731 6681 2743 6684
rect 2685 6675 2743 6681
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 6362 6672 6368 6724
rect 6420 6712 6426 6724
rect 6748 6712 6776 6740
rect 6420 6684 6776 6712
rect 6420 6672 6426 6684
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7558 6712 7564 6724
rect 7248 6684 7564 6712
rect 7248 6672 7254 6684
rect 7558 6672 7564 6684
rect 7616 6712 7622 6724
rect 8128 6712 8156 6743
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9585 6783 9643 6789
rect 8812 6774 9352 6780
rect 9585 6774 9597 6783
rect 8812 6752 9597 6774
rect 8812 6740 8818 6752
rect 9324 6749 9597 6752
rect 9631 6749 9643 6783
rect 9324 6746 9643 6749
rect 9585 6743 9643 6746
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9732 6752 10057 6780
rect 9732 6740 9738 6752
rect 10045 6749 10057 6752
rect 10091 6780 10103 6783
rect 10134 6780 10140 6792
rect 10091 6752 10140 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 10134 6740 10140 6752
rect 10192 6780 10198 6792
rect 10502 6780 10508 6792
rect 10192 6752 10508 6780
rect 10192 6740 10198 6752
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 10744 6752 11437 6780
rect 10744 6740 10750 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 7616 6684 8156 6712
rect 7616 6672 7622 6684
rect 9766 6672 9772 6724
rect 9824 6712 9830 6724
rect 9824 6684 11008 6712
rect 9824 6672 9830 6684
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 2317 6647 2375 6653
rect 2317 6644 2329 6647
rect 2096 6616 2329 6644
rect 2096 6604 2102 6616
rect 2317 6613 2329 6616
rect 2363 6613 2375 6647
rect 2317 6607 2375 6613
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 4062 6644 4068 6656
rect 3375 6616 4068 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4706 6604 4712 6656
rect 4764 6604 4770 6656
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 7340 6616 7665 6644
rect 7340 6604 7346 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 7653 6607 7711 6613
rect 9950 6604 9956 6656
rect 10008 6604 10014 6656
rect 10980 6653 11008 6684
rect 11238 6672 11244 6724
rect 11296 6712 11302 6724
rect 11669 6715 11727 6721
rect 11669 6712 11681 6715
rect 11296 6684 11681 6712
rect 11296 6672 11302 6684
rect 11669 6681 11681 6684
rect 11715 6681 11727 6715
rect 11669 6675 11727 6681
rect 11885 6715 11943 6721
rect 11885 6681 11897 6715
rect 11931 6681 11943 6715
rect 11885 6675 11943 6681
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6613 11023 6647
rect 10965 6607 11023 6613
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11900 6644 11928 6675
rect 11204 6616 11928 6644
rect 11204 6604 11210 6616
rect 1104 6554 12328 6576
rect 1104 6502 3013 6554
rect 3065 6502 3077 6554
rect 3129 6502 3141 6554
rect 3193 6502 3205 6554
rect 3257 6502 3269 6554
rect 3321 6502 5819 6554
rect 5871 6502 5883 6554
rect 5935 6502 5947 6554
rect 5999 6502 6011 6554
rect 6063 6502 6075 6554
rect 6127 6502 8625 6554
rect 8677 6502 8689 6554
rect 8741 6502 8753 6554
rect 8805 6502 8817 6554
rect 8869 6502 8881 6554
rect 8933 6502 11431 6554
rect 11483 6502 11495 6554
rect 11547 6502 11559 6554
rect 11611 6502 11623 6554
rect 11675 6502 11687 6554
rect 11739 6502 12328 6554
rect 1104 6480 12328 6502
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 3970 6440 3976 6452
rect 3927 6412 3976 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 8352 6412 8493 6440
rect 8352 6400 8358 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10686 6440 10692 6452
rect 10643 6412 10692 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 11146 6440 11152 6452
rect 10980 6412 11152 6440
rect 10980 6381 11008 6412
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11238 6400 11244 6452
rect 11296 6400 11302 6452
rect 4157 6375 4215 6381
rect 4157 6372 4169 6375
rect 3634 6344 4169 6372
rect 4157 6341 4169 6344
rect 4203 6341 4215 6375
rect 10321 6375 10379 6381
rect 10321 6372 10333 6375
rect 4157 6335 4215 6341
rect 8680 6344 10333 6372
rect 8680 6316 8708 6344
rect 10321 6341 10333 6344
rect 10367 6341 10379 6375
rect 10321 6335 10379 6341
rect 10505 6375 10563 6381
rect 10505 6341 10517 6375
rect 10551 6372 10563 6375
rect 10965 6375 11023 6381
rect 10965 6372 10977 6375
rect 10551 6344 10977 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 10965 6341 10977 6344
rect 11011 6341 11023 6375
rect 11256 6372 11284 6400
rect 10965 6335 11023 6341
rect 11072 6344 11284 6372
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 4120 6276 4261 6304
rect 4120 6264 4126 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 10100 6276 10149 6304
rect 10100 6264 10106 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6236 2191 6239
rect 2409 6239 2467 6245
rect 2179 6208 2268 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 1394 6128 1400 6180
rect 1452 6168 1458 6180
rect 2240 6168 2268 6208
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2866 6236 2872 6248
rect 2455 6208 2872 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 4154 6196 4160 6248
rect 4212 6196 4218 6248
rect 10336 6236 10364 6335
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10744 6276 10793 6304
rect 10744 6264 10750 6276
rect 10781 6273 10793 6276
rect 10827 6304 10839 6307
rect 10870 6304 10876 6316
rect 10827 6276 10876 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 11072 6313 11100 6344
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 11164 6236 11192 6267
rect 11330 6264 11336 6316
rect 11388 6264 11394 6316
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 10336 6208 11192 6236
rect 4172 6168 4200 6196
rect 1452 6140 2268 6168
rect 1452 6128 1458 6140
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1728 6072 1869 6100
rect 1728 6060 1734 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 2240 6100 2268 6140
rect 3804 6140 4200 6168
rect 3804 6100 3832 6140
rect 2240 6072 3832 6100
rect 11164 6100 11192 6208
rect 11716 6100 11744 6267
rect 11882 6128 11888 6180
rect 11940 6128 11946 6180
rect 11164 6072 11744 6100
rect 1857 6063 1915 6069
rect 1104 6010 12328 6032
rect 1104 5958 2353 6010
rect 2405 5958 2417 6010
rect 2469 5958 2481 6010
rect 2533 5958 2545 6010
rect 2597 5958 2609 6010
rect 2661 5958 5159 6010
rect 5211 5958 5223 6010
rect 5275 5958 5287 6010
rect 5339 5958 5351 6010
rect 5403 5958 5415 6010
rect 5467 5958 7965 6010
rect 8017 5958 8029 6010
rect 8081 5958 8093 6010
rect 8145 5958 8157 6010
rect 8209 5958 8221 6010
rect 8273 5958 10771 6010
rect 10823 5958 10835 6010
rect 10887 5958 10899 6010
rect 10951 5958 10963 6010
rect 11015 5958 11027 6010
rect 11079 5958 12328 6010
rect 1104 5936 12328 5958
rect 2866 5856 2872 5908
rect 2924 5856 2930 5908
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 8386 5896 8392 5908
rect 3016 5868 8392 5896
rect 3016 5856 3022 5868
rect 6380 5837 6408 5868
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8720 5868 8769 5896
rect 8720 5856 8726 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 8757 5859 8815 5865
rect 10686 5856 10692 5908
rect 10744 5856 10750 5908
rect 11793 5899 11851 5905
rect 11793 5865 11805 5899
rect 11839 5865 11851 5899
rect 11793 5859 11851 5865
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 4249 5831 4307 5837
rect 2823 5800 3464 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 1394 5720 1400 5772
rect 1452 5720 1458 5772
rect 3436 5769 3464 5800
rect 4249 5797 4261 5831
rect 4295 5797 4307 5831
rect 4249 5791 4307 5797
rect 6365 5831 6423 5837
rect 6365 5797 6377 5831
rect 6411 5797 6423 5831
rect 6365 5791 6423 5797
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5729 3479 5763
rect 3421 5723 3479 5729
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4264 5760 4292 5791
rect 10042 5788 10048 5840
rect 10100 5828 10106 5840
rect 11330 5828 11336 5840
rect 10100 5800 11336 5828
rect 10100 5788 10106 5800
rect 11330 5788 11336 5800
rect 11388 5828 11394 5840
rect 11808 5828 11836 5859
rect 11388 5800 11836 5828
rect 11388 5788 11394 5800
rect 4212 5732 7052 5760
rect 4212 5720 4218 5732
rect 7024 5704 7052 5732
rect 7282 5720 7288 5772
rect 7340 5720 7346 5772
rect 1670 5701 1676 5704
rect 1664 5692 1676 5701
rect 1631 5664 1676 5692
rect 1664 5655 1676 5664
rect 1670 5652 1676 5655
rect 1728 5652 1734 5704
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5684 5664 5917 5692
rect 5684 5652 5690 5664
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 10560 5664 10609 5692
rect 10560 5652 10566 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 10686 5652 10692 5704
rect 10744 5692 10750 5704
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 10744 5664 10793 5692
rect 10744 5652 10750 5664
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 5813 5627 5871 5633
rect 5813 5624 5825 5627
rect 4580 5596 5825 5624
rect 4580 5584 4586 5596
rect 5813 5593 5825 5596
rect 5859 5624 5871 5627
rect 6178 5624 6184 5636
rect 5859 5596 6184 5624
rect 5859 5593 5871 5596
rect 5813 5587 5871 5593
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 6362 5584 6368 5636
rect 6420 5584 6426 5636
rect 8294 5584 8300 5636
rect 8352 5584 8358 5636
rect 5626 5516 5632 5568
rect 5684 5516 5690 5568
rect 1104 5466 12328 5488
rect 1104 5414 3013 5466
rect 3065 5414 3077 5466
rect 3129 5414 3141 5466
rect 3193 5414 3205 5466
rect 3257 5414 3269 5466
rect 3321 5414 5819 5466
rect 5871 5414 5883 5466
rect 5935 5414 5947 5466
rect 5999 5414 6011 5466
rect 6063 5414 6075 5466
rect 6127 5414 8625 5466
rect 8677 5414 8689 5466
rect 8741 5414 8753 5466
rect 8805 5414 8817 5466
rect 8869 5414 8881 5466
rect 8933 5414 11431 5466
rect 11483 5414 11495 5466
rect 11547 5414 11559 5466
rect 11611 5414 11623 5466
rect 11675 5414 11687 5466
rect 11739 5414 12328 5466
rect 1104 5392 12328 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4120 5324 5672 5352
rect 4120 5312 4126 5324
rect 4614 5244 4620 5296
rect 4672 5244 4678 5296
rect 5644 5284 5672 5324
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5776 5324 5825 5352
rect 5776 5312 5782 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 6362 5312 6368 5364
rect 6420 5312 6426 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8294 5352 8300 5364
rect 7975 5324 8300 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 7742 5284 7748 5296
rect 5644 5256 7748 5284
rect 7742 5244 7748 5256
rect 7800 5284 7806 5296
rect 7800 5256 7880 5284
rect 7800 5244 7806 5256
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6227 5188 6561 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6549 5185 6561 5188
rect 6595 5216 6607 5219
rect 6914 5216 6920 5228
rect 6595 5188 6920 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 3743 5120 3832 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 3804 5012 3832 5120
rect 3970 5108 3976 5160
rect 4028 5108 4034 5160
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 6012 5148 6040 5179
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7852 5225 7880 5256
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 11974 5176 11980 5228
rect 12032 5176 12038 5228
rect 6733 5151 6791 5157
rect 6733 5148 6745 5151
rect 5776 5120 6745 5148
rect 5776 5108 5782 5120
rect 6733 5117 6745 5120
rect 6779 5148 6791 5151
rect 7374 5148 7380 5160
rect 6779 5120 7380 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 7374 5108 7380 5120
rect 7432 5148 7438 5160
rect 10502 5148 10508 5160
rect 7432 5120 10508 5148
rect 7432 5108 7438 5120
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 4154 5012 4160 5024
rect 3804 4984 4160 5012
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 10744 4984 11805 5012
rect 10744 4972 10750 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 11793 4975 11851 4981
rect 1104 4922 12328 4944
rect 1104 4870 2353 4922
rect 2405 4870 2417 4922
rect 2469 4870 2481 4922
rect 2533 4870 2545 4922
rect 2597 4870 2609 4922
rect 2661 4870 5159 4922
rect 5211 4870 5223 4922
rect 5275 4870 5287 4922
rect 5339 4870 5351 4922
rect 5403 4870 5415 4922
rect 5467 4870 7965 4922
rect 8017 4870 8029 4922
rect 8081 4870 8093 4922
rect 8145 4870 8157 4922
rect 8209 4870 8221 4922
rect 8273 4870 10771 4922
rect 10823 4870 10835 4922
rect 10887 4870 10899 4922
rect 10951 4870 10963 4922
rect 11015 4870 11027 4922
rect 11079 4870 12328 4922
rect 1104 4848 12328 4870
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4801 4811 4859 4817
rect 4801 4808 4813 4811
rect 4028 4780 4813 4808
rect 4028 4768 4034 4780
rect 4801 4777 4813 4780
rect 4847 4777 4859 4811
rect 5534 4808 5540 4820
rect 4801 4771 4859 4777
rect 5276 4780 5540 4808
rect 4614 4700 4620 4752
rect 4672 4700 4678 4752
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4120 4576 4537 4604
rect 4120 4564 4126 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4764 4576 4997 4604
rect 4764 4564 4770 4576
rect 4985 4573 4997 4576
rect 5031 4604 5043 4607
rect 5276 4604 5304 4780
rect 5534 4768 5540 4780
rect 5592 4808 5598 4820
rect 9030 4808 9036 4820
rect 5592 4780 9036 4808
rect 5592 4768 5598 4780
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9640 4780 9873 4808
rect 9640 4768 9646 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 9861 4771 9919 4777
rect 10321 4811 10379 4817
rect 10321 4777 10333 4811
rect 10367 4777 10379 4811
rect 10321 4771 10379 4777
rect 8386 4700 8392 4752
rect 8444 4740 8450 4752
rect 8941 4743 8999 4749
rect 8941 4740 8953 4743
rect 8444 4712 8953 4740
rect 8444 4700 8450 4712
rect 8941 4709 8953 4712
rect 8987 4709 8999 4743
rect 10336 4740 10364 4771
rect 10686 4740 10692 4752
rect 10336 4712 10692 4740
rect 8941 4703 8999 4709
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 9493 4675 9551 4681
rect 9493 4672 9505 4675
rect 5368 4644 9505 4672
rect 5368 4613 5396 4644
rect 9493 4641 9505 4644
rect 9539 4641 9551 4675
rect 9493 4635 9551 4641
rect 10226 4632 10232 4684
rect 10284 4632 10290 4684
rect 5031 4576 5304 4604
rect 5353 4607 5411 4613
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5626 4604 5632 4616
rect 5491 4576 5632 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 9088 4576 9137 4604
rect 9088 4564 9094 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 10502 4564 10508 4616
rect 10560 4564 10566 4616
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 3878 4496 3884 4548
rect 3936 4536 3942 4548
rect 5077 4539 5135 4545
rect 5077 4536 5089 4539
rect 3936 4508 5089 4536
rect 3936 4496 3942 4508
rect 5077 4505 5089 4508
rect 5123 4505 5135 4539
rect 5077 4499 5135 4505
rect 5169 4539 5227 4545
rect 5169 4505 5181 4539
rect 5215 4536 5227 4539
rect 5718 4536 5724 4548
rect 5215 4508 5724 4536
rect 5215 4505 5227 4508
rect 5169 4499 5227 4505
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 7558 4536 7564 4548
rect 6972 4508 7564 4536
rect 6972 4496 6978 4508
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 9217 4539 9275 4545
rect 9217 4505 9229 4539
rect 9263 4536 9275 4539
rect 10134 4536 10140 4548
rect 9263 4508 10140 4536
rect 9263 4505 9275 4508
rect 9217 4499 9275 4505
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 10321 4539 10379 4545
rect 10321 4505 10333 4539
rect 10367 4505 10379 4539
rect 10321 4499 10379 4505
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 8294 4468 8300 4480
rect 6236 4440 8300 4468
rect 6236 4428 6242 4440
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 9306 4428 9312 4480
rect 9364 4428 9370 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10336 4468 10364 4499
rect 11238 4496 11244 4548
rect 11296 4496 11302 4548
rect 9732 4440 10364 4468
rect 9732 4428 9738 4440
rect 1104 4378 12328 4400
rect 1104 4326 3013 4378
rect 3065 4326 3077 4378
rect 3129 4326 3141 4378
rect 3193 4326 3205 4378
rect 3257 4326 3269 4378
rect 3321 4326 5819 4378
rect 5871 4326 5883 4378
rect 5935 4326 5947 4378
rect 5999 4326 6011 4378
rect 6063 4326 6075 4378
rect 6127 4326 8625 4378
rect 8677 4326 8689 4378
rect 8741 4326 8753 4378
rect 8805 4326 8817 4378
rect 8869 4326 8881 4378
rect 8933 4326 11431 4378
rect 11483 4326 11495 4378
rect 11547 4326 11559 4378
rect 11611 4326 11623 4378
rect 11675 4326 11687 4378
rect 11739 4326 12328 4378
rect 1104 4304 12328 4326
rect 2777 4267 2835 4273
rect 2777 4233 2789 4267
rect 2823 4264 2835 4267
rect 4706 4264 4712 4276
rect 2823 4236 4712 4264
rect 2823 4233 2835 4236
rect 2777 4227 2835 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8444 4236 8493 4264
rect 8444 4224 8450 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 9364 4236 9597 4264
rect 9364 4224 9370 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 9585 4227 9643 4233
rect 9876 4236 11652 4264
rect 6822 4196 6828 4208
rect 6564 4168 6828 4196
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2188 4100 2697 4128
rect 2188 4088 2194 4100
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3016 4100 3893 4128
rect 3016 4088 3022 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 6178 4128 6184 4140
rect 5583 4100 6184 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 2884 3992 2912 4023
rect 3602 4020 3608 4072
rect 3660 4020 3666 4072
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 6564 4060 6592 4168
rect 6822 4156 6828 4168
rect 6880 4196 6886 4208
rect 8113 4199 8171 4205
rect 6880 4168 7420 4196
rect 6880 4156 6886 4168
rect 6914 4088 6920 4140
rect 6972 4088 6978 4140
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 5859 4032 6592 4060
rect 7116 4060 7144 4091
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 7392 4137 7420 4168
rect 8113 4165 8125 4199
rect 8159 4196 8171 4199
rect 9030 4196 9036 4208
rect 8159 4168 9036 4196
rect 8159 4165 8171 4168
rect 8113 4159 8171 4165
rect 9030 4156 9036 4168
rect 9088 4196 9094 4208
rect 9876 4196 9904 4236
rect 9088 4168 9904 4196
rect 9088 4156 9094 4168
rect 10226 4156 10232 4208
rect 10284 4196 10290 4208
rect 10284 4168 10640 4196
rect 10284 4156 10290 4168
rect 10612 4140 10640 4168
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7650 4088 7656 4140
rect 7708 4088 7714 4140
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 8938 4128 8944 4140
rect 8619 4100 8944 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9766 4088 9772 4140
rect 9824 4088 9830 4140
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 10091 4100 10548 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 7834 4060 7840 4072
rect 7116 4032 7840 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 7834 4020 7840 4032
rect 7892 4060 7898 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7892 4032 7941 4060
rect 7892 4020 7898 4032
rect 7929 4029 7941 4032
rect 7975 4060 7987 4063
rect 10410 4060 10416 4072
rect 7975 4032 10416 4060
rect 7975 4029 7987 4032
rect 7929 4023 7987 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 10520 4060 10548 4100
rect 10594 4088 10600 4140
rect 10652 4088 10658 4140
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11238 4128 11244 4140
rect 11195 4100 11244 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11238 4088 11244 4100
rect 11296 4128 11302 4140
rect 11624 4137 11652 4236
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11296 4100 11529 4128
rect 11296 4088 11302 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 10520 4032 11192 4060
rect 2740 3964 2912 3992
rect 5629 3995 5687 4001
rect 2740 3952 2746 3964
rect 5629 3961 5641 3995
rect 5675 3992 5687 3995
rect 6086 3992 6092 4004
rect 5675 3964 6092 3992
rect 5675 3961 5687 3964
rect 5629 3955 5687 3961
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 7558 3952 7564 4004
rect 7616 3992 7622 4004
rect 8297 3995 8355 4001
rect 8297 3992 8309 3995
rect 7616 3964 8309 3992
rect 7616 3952 7622 3964
rect 8297 3961 8309 3964
rect 8343 3961 8355 3995
rect 8297 3955 8355 3961
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 10226 3992 10232 4004
rect 10008 3964 10232 3992
rect 10008 3952 10014 3964
rect 10226 3952 10232 3964
rect 10284 3992 10290 4004
rect 11057 3995 11115 4001
rect 11057 3992 11069 3995
rect 10284 3964 11069 3992
rect 10284 3952 10290 3964
rect 11057 3961 11069 3964
rect 11103 3961 11115 3995
rect 11164 3992 11192 4032
rect 11164 3964 11652 3992
rect 11057 3955 11115 3961
rect 11624 3936 11652 3964
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 2317 3927 2375 3933
rect 2317 3924 2329 3927
rect 1820 3896 2329 3924
rect 1820 3884 1826 3896
rect 2317 3893 2329 3896
rect 2363 3893 2375 3927
rect 2317 3887 2375 3893
rect 5721 3927 5779 3933
rect 5721 3893 5733 3927
rect 5767 3924 5779 3927
rect 6454 3924 6460 3936
rect 5767 3896 6460 3924
rect 5767 3893 5779 3896
rect 5721 3887 5779 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 7377 3927 7435 3933
rect 7377 3893 7389 3927
rect 7423 3924 7435 3927
rect 7466 3924 7472 3936
rect 7423 3896 7472 3924
rect 7423 3893 7435 3896
rect 7377 3887 7435 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 10652 3896 11529 3924
rect 10652 3884 10658 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 11664 3896 11897 3924
rect 11664 3884 11670 3896
rect 11885 3893 11897 3896
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 1104 3834 12328 3856
rect 1104 3782 2353 3834
rect 2405 3782 2417 3834
rect 2469 3782 2481 3834
rect 2533 3782 2545 3834
rect 2597 3782 2609 3834
rect 2661 3782 5159 3834
rect 5211 3782 5223 3834
rect 5275 3782 5287 3834
rect 5339 3782 5351 3834
rect 5403 3782 5415 3834
rect 5467 3782 7965 3834
rect 8017 3782 8029 3834
rect 8081 3782 8093 3834
rect 8145 3782 8157 3834
rect 8209 3782 8221 3834
rect 8273 3782 10771 3834
rect 10823 3782 10835 3834
rect 10887 3782 10899 3834
rect 10951 3782 10963 3834
rect 11015 3782 11027 3834
rect 11079 3782 12328 3834
rect 1104 3760 12328 3782
rect 3602 3680 3608 3732
rect 3660 3680 3666 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3936 3692 3985 3720
rect 3936 3680 3942 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 6914 3720 6920 3732
rect 3973 3683 4031 3689
rect 6564 3692 6920 3720
rect 3988 3652 4016 3683
rect 3988 3624 5948 3652
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 1452 3556 1869 3584
rect 1452 3544 1458 3556
rect 1857 3553 1869 3556
rect 1903 3584 1915 3587
rect 4154 3584 4160 3596
rect 1903 3556 4160 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 1762 3476 1768 3528
rect 1820 3476 1826 3528
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3660 3488 3893 3516
rect 3660 3476 3666 3488
rect 3881 3485 3893 3488
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 5626 3516 5632 3528
rect 5583 3488 5632 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 5920 3525 5948 3624
rect 6454 3544 6460 3596
rect 6512 3544 6518 3596
rect 6564 3593 6592 3692
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 7650 3720 7656 3732
rect 7147 3692 7656 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 7926 3720 7932 3732
rect 7791 3692 7932 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 8938 3680 8944 3732
rect 8996 3680 9002 3732
rect 9585 3723 9643 3729
rect 9585 3689 9597 3723
rect 9631 3720 9643 3723
rect 9674 3720 9680 3732
rect 9631 3692 9680 3720
rect 9631 3689 9643 3692
rect 9585 3683 9643 3689
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10134 3680 10140 3732
rect 10192 3680 10198 3732
rect 8665 3655 8723 3661
rect 8665 3652 8677 3655
rect 6656 3624 8677 3652
rect 6656 3593 6684 3624
rect 8665 3621 8677 3624
rect 8711 3621 8723 3655
rect 8665 3615 8723 3621
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 6641 3587 6699 3593
rect 6641 3553 6653 3587
rect 6687 3553 6699 3587
rect 7282 3584 7288 3596
rect 6641 3547 6699 3553
rect 7024 3556 7288 3584
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 2130 3408 2136 3460
rect 2188 3408 2194 3460
rect 3694 3448 3700 3460
rect 3358 3420 3700 3448
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 5828 3448 5856 3479
rect 6086 3448 6092 3460
rect 5828 3420 6092 3448
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 6181 3451 6239 3457
rect 6181 3417 6193 3451
rect 6227 3448 6239 3451
rect 6748 3448 6776 3479
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 7024 3525 7052 3556
rect 7282 3544 7288 3556
rect 7340 3584 7346 3596
rect 7340 3556 8616 3584
rect 7340 3544 7346 3556
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6880 3488 7021 3516
rect 6880 3476 6886 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 6227 3420 6776 3448
rect 7208 3448 7236 3479
rect 7466 3476 7472 3528
rect 7524 3476 7530 3528
rect 7558 3476 7564 3528
rect 7616 3476 7622 3528
rect 7834 3476 7840 3528
rect 7892 3476 7898 3528
rect 8588 3525 8616 3556
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 7852 3448 7880 3476
rect 7208 3420 7880 3448
rect 6227 3417 6239 3420
rect 6181 3411 6239 3417
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 1670 3380 1676 3392
rect 1627 3352 1676 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 6270 3340 6276 3392
rect 6328 3340 6334 3392
rect 7282 3340 7288 3392
rect 7340 3340 7346 3392
rect 7742 3340 7748 3392
rect 7800 3380 7806 3392
rect 7944 3380 7972 3479
rect 7800 3352 7972 3380
rect 7800 3340 7806 3352
rect 8018 3340 8024 3392
rect 8076 3340 8082 3392
rect 8588 3380 8616 3479
rect 8680 3448 8708 3615
rect 9766 3612 9772 3664
rect 9824 3612 9830 3664
rect 10594 3612 10600 3664
rect 10652 3652 10658 3664
rect 11701 3655 11759 3661
rect 11701 3652 11713 3655
rect 10652 3624 11713 3652
rect 10652 3612 10658 3624
rect 11701 3621 11713 3624
rect 11747 3621 11759 3655
rect 11701 3615 11759 3621
rect 9784 3584 9812 3612
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9140 3556 9965 3584
rect 9140 3525 9168 3556
rect 9953 3553 9965 3556
rect 9999 3584 10011 3587
rect 9999 3556 10088 3584
rect 9999 3553 10011 3556
rect 9953 3547 10011 3553
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9398 3476 9404 3528
rect 9456 3476 9462 3528
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 8680 3420 9321 3448
rect 9309 3417 9321 3420
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 9508 3380 9536 3479
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 10060 3525 10088 3556
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3516 10747 3519
rect 11606 3516 11612 3528
rect 10735 3488 11612 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 11882 3408 11888 3460
rect 11940 3408 11946 3460
rect 8588 3352 9536 3380
rect 1104 3290 12328 3312
rect 1104 3238 3013 3290
rect 3065 3238 3077 3290
rect 3129 3238 3141 3290
rect 3193 3238 3205 3290
rect 3257 3238 3269 3290
rect 3321 3238 5819 3290
rect 5871 3238 5883 3290
rect 5935 3238 5947 3290
rect 5999 3238 6011 3290
rect 6063 3238 6075 3290
rect 6127 3238 8625 3290
rect 8677 3238 8689 3290
rect 8741 3238 8753 3290
rect 8805 3238 8817 3290
rect 8869 3238 8881 3290
rect 8933 3238 11431 3290
rect 11483 3238 11495 3290
rect 11547 3238 11559 3290
rect 11611 3238 11623 3290
rect 11675 3238 11687 3290
rect 11739 3238 12328 3290
rect 1104 3216 12328 3238
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 2869 3179 2927 3185
rect 2869 3176 2881 3179
rect 2188 3148 2881 3176
rect 2188 3136 2194 3148
rect 2869 3145 2881 3148
rect 2915 3145 2927 3179
rect 2869 3139 2927 3145
rect 3694 3136 3700 3188
rect 3752 3136 3758 3188
rect 6270 3176 6276 3188
rect 4448 3148 6276 3176
rect 4448 3117 4476 3148
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7190 3176 7196 3188
rect 6972 3148 7196 3176
rect 6972 3136 6978 3148
rect 7190 3136 7196 3148
rect 7248 3176 7254 3188
rect 7926 3176 7932 3188
rect 7248 3148 7932 3176
rect 7248 3136 7254 3148
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9030 3176 9036 3188
rect 8803 3148 9036 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9456 3148 9873 3176
rect 9456 3136 9462 3148
rect 9861 3145 9873 3148
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 4433 3111 4491 3117
rect 4433 3077 4445 3111
rect 4479 3077 4491 3111
rect 4433 3071 4491 3077
rect 7282 3068 7288 3120
rect 7340 3068 7346 3120
rect 8018 3068 8024 3120
rect 8076 3068 8082 3120
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 9732 3080 9996 3108
rect 9732 3068 9738 3080
rect 1394 3000 1400 3052
rect 1452 3000 1458 3052
rect 1670 3049 1676 3052
rect 1664 3040 1676 3049
rect 1631 3012 1676 3040
rect 1664 3003 1676 3012
rect 1670 3000 1676 3003
rect 1728 3000 1734 3052
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4062 3040 4068 3052
rect 3835 3012 4068 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4154 3000 4160 3052
rect 4212 3000 4218 3052
rect 5534 3000 5540 3052
rect 5592 3000 5598 3052
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 9968 3049 9996 3080
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10468 3012 10701 3040
rect 10468 3000 10474 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 2777 2907 2835 2913
rect 2777 2873 2789 2907
rect 2823 2904 2835 2907
rect 3436 2904 3464 2935
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 5905 2975 5963 2981
rect 5905 2972 5917 2975
rect 5684 2944 5917 2972
rect 5684 2932 5690 2944
rect 5905 2941 5917 2944
rect 5951 2972 5963 2975
rect 6822 2972 6828 2984
rect 5951 2944 6828 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 9784 2972 9812 3000
rect 9784 2944 10364 2972
rect 10336 2913 10364 2944
rect 10594 2932 10600 2984
rect 10652 2932 10658 2984
rect 2823 2876 3464 2904
rect 10321 2907 10379 2913
rect 2823 2873 2835 2876
rect 2777 2867 2835 2873
rect 10321 2873 10333 2907
rect 10367 2873 10379 2907
rect 10321 2867 10379 2873
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 9674 2836 9680 2848
rect 6236 2808 9680 2836
rect 6236 2796 6242 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 1104 2746 12328 2768
rect 1104 2694 2353 2746
rect 2405 2694 2417 2746
rect 2469 2694 2481 2746
rect 2533 2694 2545 2746
rect 2597 2694 2609 2746
rect 2661 2694 5159 2746
rect 5211 2694 5223 2746
rect 5275 2694 5287 2746
rect 5339 2694 5351 2746
rect 5403 2694 5415 2746
rect 5467 2694 7965 2746
rect 8017 2694 8029 2746
rect 8081 2694 8093 2746
rect 8145 2694 8157 2746
rect 8209 2694 8221 2746
rect 8273 2694 10771 2746
rect 10823 2694 10835 2746
rect 10887 2694 10899 2746
rect 10951 2694 10963 2746
rect 11015 2694 11027 2746
rect 11079 2694 12328 2746
rect 1104 2672 12328 2694
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5534 2632 5540 2644
rect 5215 2604 5540 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6178 2632 6184 2644
rect 6135 2604 6184 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 7432 2468 8156 2496
rect 7432 2456 7438 2468
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 4120 2400 5089 2428
rect 4120 2388 4126 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5776 2400 5917 2428
rect 5776 2388 5782 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6822 2388 6828 2440
rect 6880 2388 6886 2440
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7650 2428 7656 2440
rect 7515 2400 7656 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8128 2437 8156 2468
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7156 2264 7297 2292
rect 7156 2252 7162 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7800 2264 7941 2292
rect 7800 2252 7806 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 1104 2202 12328 2224
rect 1104 2150 3013 2202
rect 3065 2150 3077 2202
rect 3129 2150 3141 2202
rect 3193 2150 3205 2202
rect 3257 2150 3269 2202
rect 3321 2150 5819 2202
rect 5871 2150 5883 2202
rect 5935 2150 5947 2202
rect 5999 2150 6011 2202
rect 6063 2150 6075 2202
rect 6127 2150 8625 2202
rect 8677 2150 8689 2202
rect 8741 2150 8753 2202
rect 8805 2150 8817 2202
rect 8869 2150 8881 2202
rect 8933 2150 11431 2202
rect 11483 2150 11495 2202
rect 11547 2150 11559 2202
rect 11611 2150 11623 2202
rect 11675 2150 11687 2202
rect 11739 2150 12328 2202
rect 1104 2128 12328 2150
<< via1 >>
rect 3013 13030 3065 13082
rect 3077 13030 3129 13082
rect 3141 13030 3193 13082
rect 3205 13030 3257 13082
rect 3269 13030 3321 13082
rect 5819 13030 5871 13082
rect 5883 13030 5935 13082
rect 5947 13030 5999 13082
rect 6011 13030 6063 13082
rect 6075 13030 6127 13082
rect 8625 13030 8677 13082
rect 8689 13030 8741 13082
rect 8753 13030 8805 13082
rect 8817 13030 8869 13082
rect 8881 13030 8933 13082
rect 11431 13030 11483 13082
rect 11495 13030 11547 13082
rect 11559 13030 11611 13082
rect 11623 13030 11675 13082
rect 11687 13030 11739 13082
rect 5724 12928 5776 12980
rect 6460 12860 6512 12912
rect 5540 12792 5592 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7104 12792 7156 12844
rect 7748 12792 7800 12844
rect 8392 12792 8444 12844
rect 7564 12588 7616 12640
rect 8300 12588 8352 12640
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 2353 12486 2405 12538
rect 2417 12486 2469 12538
rect 2481 12486 2533 12538
rect 2545 12486 2597 12538
rect 2609 12486 2661 12538
rect 5159 12486 5211 12538
rect 5223 12486 5275 12538
rect 5287 12486 5339 12538
rect 5351 12486 5403 12538
rect 5415 12486 5467 12538
rect 7965 12486 8017 12538
rect 8029 12486 8081 12538
rect 8093 12486 8145 12538
rect 8157 12486 8209 12538
rect 8221 12486 8273 12538
rect 10771 12486 10823 12538
rect 10835 12486 10887 12538
rect 10899 12486 10951 12538
rect 10963 12486 11015 12538
rect 11027 12486 11079 12538
rect 6184 12316 6236 12368
rect 2596 12248 2648 12300
rect 4988 12180 5040 12232
rect 1584 12155 1636 12164
rect 1584 12121 1593 12155
rect 1593 12121 1627 12155
rect 1627 12121 1636 12155
rect 1584 12112 1636 12121
rect 2320 12112 2372 12164
rect 4528 12112 4580 12164
rect 5540 12112 5592 12164
rect 7380 12223 7432 12232
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 7564 12112 7616 12164
rect 8300 12180 8352 12232
rect 10324 12180 10376 12232
rect 11244 12180 11296 12232
rect 5632 12044 5684 12096
rect 8392 12112 8444 12164
rect 9864 12155 9916 12164
rect 9864 12121 9873 12155
rect 9873 12121 9907 12155
rect 9907 12121 9916 12155
rect 9864 12112 9916 12121
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 8116 12044 8168 12096
rect 9312 12044 9364 12096
rect 3013 11942 3065 11994
rect 3077 11942 3129 11994
rect 3141 11942 3193 11994
rect 3205 11942 3257 11994
rect 3269 11942 3321 11994
rect 5819 11942 5871 11994
rect 5883 11942 5935 11994
rect 5947 11942 5999 11994
rect 6011 11942 6063 11994
rect 6075 11942 6127 11994
rect 8625 11942 8677 11994
rect 8689 11942 8741 11994
rect 8753 11942 8805 11994
rect 8817 11942 8869 11994
rect 8881 11942 8933 11994
rect 11431 11942 11483 11994
rect 11495 11942 11547 11994
rect 11559 11942 11611 11994
rect 11623 11942 11675 11994
rect 11687 11942 11739 11994
rect 2320 11840 2372 11892
rect 5540 11840 5592 11892
rect 7380 11840 7432 11892
rect 2780 11772 2832 11824
rect 3332 11772 3384 11824
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 4896 11704 4948 11756
rect 5540 11704 5592 11756
rect 6184 11772 6236 11824
rect 7932 11772 7984 11824
rect 6368 11704 6420 11756
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 7748 11704 7800 11756
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 8392 11704 8444 11756
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 6184 11568 6236 11620
rect 6644 11568 6696 11620
rect 8116 11679 8168 11688
rect 8116 11645 8125 11679
rect 8125 11645 8159 11679
rect 8159 11645 8168 11679
rect 8116 11636 8168 11645
rect 9864 11636 9916 11688
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 10692 11704 10744 11756
rect 11152 11704 11204 11756
rect 11336 11636 11388 11688
rect 4712 11500 4764 11552
rect 8392 11568 8444 11620
rect 2353 11398 2405 11450
rect 2417 11398 2469 11450
rect 2481 11398 2533 11450
rect 2545 11398 2597 11450
rect 2609 11398 2661 11450
rect 5159 11398 5211 11450
rect 5223 11398 5275 11450
rect 5287 11398 5339 11450
rect 5351 11398 5403 11450
rect 5415 11398 5467 11450
rect 7965 11398 8017 11450
rect 8029 11398 8081 11450
rect 8093 11398 8145 11450
rect 8157 11398 8209 11450
rect 8221 11398 8273 11450
rect 10771 11398 10823 11450
rect 10835 11398 10887 11450
rect 10899 11398 10951 11450
rect 10963 11398 11015 11450
rect 11027 11398 11079 11450
rect 3332 11296 3384 11348
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 4896 11339 4948 11348
rect 4896 11305 4905 11339
rect 4905 11305 4939 11339
rect 4939 11305 4948 11339
rect 4896 11296 4948 11305
rect 2780 11228 2832 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 7012 11296 7064 11348
rect 7472 11296 7524 11348
rect 8392 11296 8444 11348
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 11336 11228 11388 11280
rect 3424 11092 3476 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 7656 11160 7708 11212
rect 1584 11024 1636 11076
rect 4988 11024 5040 11076
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6552 11092 6604 11144
rect 6644 11092 6696 11144
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 11152 11092 11204 11101
rect 7380 11024 7432 11076
rect 8392 11024 8444 11076
rect 5356 10999 5408 11008
rect 5356 10965 5365 10999
rect 5365 10965 5399 10999
rect 5399 10965 5408 10999
rect 5356 10956 5408 10965
rect 3013 10854 3065 10906
rect 3077 10854 3129 10906
rect 3141 10854 3193 10906
rect 3205 10854 3257 10906
rect 3269 10854 3321 10906
rect 5819 10854 5871 10906
rect 5883 10854 5935 10906
rect 5947 10854 5999 10906
rect 6011 10854 6063 10906
rect 6075 10854 6127 10906
rect 8625 10854 8677 10906
rect 8689 10854 8741 10906
rect 8753 10854 8805 10906
rect 8817 10854 8869 10906
rect 8881 10854 8933 10906
rect 11431 10854 11483 10906
rect 11495 10854 11547 10906
rect 11559 10854 11611 10906
rect 11623 10854 11675 10906
rect 11687 10854 11739 10906
rect 5356 10752 5408 10804
rect 6368 10795 6420 10804
rect 6368 10761 6377 10795
rect 6377 10761 6411 10795
rect 6411 10761 6420 10795
rect 6368 10752 6420 10761
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 6920 10684 6972 10736
rect 8484 10727 8536 10736
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 7564 10616 7616 10668
rect 8484 10693 8493 10727
rect 8493 10693 8527 10727
rect 8527 10693 8536 10727
rect 8484 10684 8536 10693
rect 10692 10752 10744 10804
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 10416 10684 10468 10736
rect 8576 10616 8628 10668
rect 9864 10616 9916 10668
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11152 10616 11204 10668
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 10140 10548 10192 10600
rect 10876 10548 10928 10600
rect 5724 10480 5776 10532
rect 5908 10480 5960 10532
rect 9588 10480 9640 10532
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 2353 10310 2405 10362
rect 2417 10310 2469 10362
rect 2481 10310 2533 10362
rect 2545 10310 2597 10362
rect 2609 10310 2661 10362
rect 5159 10310 5211 10362
rect 5223 10310 5275 10362
rect 5287 10310 5339 10362
rect 5351 10310 5403 10362
rect 5415 10310 5467 10362
rect 7965 10310 8017 10362
rect 8029 10310 8081 10362
rect 8093 10310 8145 10362
rect 8157 10310 8209 10362
rect 8221 10310 8273 10362
rect 10771 10310 10823 10362
rect 10835 10310 10887 10362
rect 10899 10310 10951 10362
rect 10963 10310 11015 10362
rect 11027 10310 11079 10362
rect 1308 10208 1360 10260
rect 5080 10208 5132 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 1584 10004 1636 10056
rect 6000 10140 6052 10192
rect 6000 10047 6052 10056
rect 5080 9936 5132 9988
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 9128 10140 9180 10192
rect 9864 10115 9916 10124
rect 9864 10081 9873 10115
rect 9873 10081 9907 10115
rect 9907 10081 9916 10115
rect 9864 10072 9916 10081
rect 8484 10004 8536 10056
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 6368 9936 6420 9988
rect 8576 9936 8628 9988
rect 9404 9979 9456 9988
rect 9404 9945 9413 9979
rect 9413 9945 9447 9979
rect 9447 9945 9456 9979
rect 9404 9936 9456 9945
rect 6460 9868 6512 9920
rect 9312 9868 9364 9920
rect 3013 9766 3065 9818
rect 3077 9766 3129 9818
rect 3141 9766 3193 9818
rect 3205 9766 3257 9818
rect 3269 9766 3321 9818
rect 5819 9766 5871 9818
rect 5883 9766 5935 9818
rect 5947 9766 5999 9818
rect 6011 9766 6063 9818
rect 6075 9766 6127 9818
rect 8625 9766 8677 9818
rect 8689 9766 8741 9818
rect 8753 9766 8805 9818
rect 8817 9766 8869 9818
rect 8881 9766 8933 9818
rect 11431 9766 11483 9818
rect 11495 9766 11547 9818
rect 11559 9766 11611 9818
rect 11623 9766 11675 9818
rect 11687 9766 11739 9818
rect 7288 9639 7340 9648
rect 7288 9605 7297 9639
rect 7297 9605 7331 9639
rect 7331 9605 7340 9639
rect 7288 9596 7340 9605
rect 9864 9664 9916 9716
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 2780 9528 2832 9580
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 6460 9528 6512 9580
rect 6828 9528 6880 9580
rect 9404 9528 9456 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 2688 9460 2740 9512
rect 6552 9460 6604 9512
rect 7472 9460 7524 9512
rect 9128 9460 9180 9512
rect 11336 9392 11388 9444
rect 2688 9324 2740 9376
rect 5540 9324 5592 9376
rect 5908 9324 5960 9376
rect 2353 9222 2405 9274
rect 2417 9222 2469 9274
rect 2481 9222 2533 9274
rect 2545 9222 2597 9274
rect 2609 9222 2661 9274
rect 5159 9222 5211 9274
rect 5223 9222 5275 9274
rect 5287 9222 5339 9274
rect 5351 9222 5403 9274
rect 5415 9222 5467 9274
rect 7965 9222 8017 9274
rect 8029 9222 8081 9274
rect 8093 9222 8145 9274
rect 8157 9222 8209 9274
rect 8221 9222 8273 9274
rect 10771 9222 10823 9274
rect 10835 9222 10887 9274
rect 10899 9222 10951 9274
rect 10963 9222 11015 9274
rect 11027 9222 11079 9274
rect 1676 9120 1728 9172
rect 2780 9120 2832 9172
rect 5908 9163 5960 9172
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 8300 9120 8352 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 10508 9120 10560 9172
rect 10692 9052 10744 9104
rect 2688 8984 2740 9036
rect 5724 9027 5776 9036
rect 5724 8993 5733 9027
rect 5733 8993 5767 9027
rect 5767 8993 5776 9027
rect 5724 8984 5776 8993
rect 7472 8984 7524 9036
rect 9404 8984 9456 9036
rect 3424 8916 3476 8968
rect 3792 8916 3844 8968
rect 4896 8916 4948 8968
rect 5264 8916 5316 8968
rect 5540 8848 5592 8900
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 7472 8891 7524 8900
rect 7472 8857 7481 8891
rect 7481 8857 7515 8891
rect 7515 8857 7524 8891
rect 7472 8848 7524 8857
rect 8300 8848 8352 8900
rect 7012 8780 7064 8832
rect 7564 8823 7616 8832
rect 7564 8789 7573 8823
rect 7573 8789 7607 8823
rect 7607 8789 7616 8823
rect 7564 8780 7616 8789
rect 8208 8823 8260 8832
rect 8208 8789 8217 8823
rect 8217 8789 8251 8823
rect 8251 8789 8260 8823
rect 8208 8780 8260 8789
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 3013 8678 3065 8730
rect 3077 8678 3129 8730
rect 3141 8678 3193 8730
rect 3205 8678 3257 8730
rect 3269 8678 3321 8730
rect 5819 8678 5871 8730
rect 5883 8678 5935 8730
rect 5947 8678 5999 8730
rect 6011 8678 6063 8730
rect 6075 8678 6127 8730
rect 8625 8678 8677 8730
rect 8689 8678 8741 8730
rect 8753 8678 8805 8730
rect 8817 8678 8869 8730
rect 8881 8678 8933 8730
rect 11431 8678 11483 8730
rect 11495 8678 11547 8730
rect 11559 8678 11611 8730
rect 11623 8678 11675 8730
rect 11687 8678 11739 8730
rect 2688 8576 2740 8628
rect 5724 8576 5776 8628
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 8208 8576 8260 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 6644 8508 6696 8560
rect 2964 8372 3016 8424
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 4160 8236 4212 8288
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 5080 8236 5132 8288
rect 5540 8304 5592 8356
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 8392 8440 8444 8492
rect 9036 8508 9088 8560
rect 11060 8508 11112 8560
rect 10048 8440 10100 8492
rect 10140 8440 10192 8492
rect 8300 8372 8352 8424
rect 10416 8372 10468 8424
rect 6552 8236 6604 8288
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 2353 8134 2405 8186
rect 2417 8134 2469 8186
rect 2481 8134 2533 8186
rect 2545 8134 2597 8186
rect 2609 8134 2661 8186
rect 5159 8134 5211 8186
rect 5223 8134 5275 8186
rect 5287 8134 5339 8186
rect 5351 8134 5403 8186
rect 5415 8134 5467 8186
rect 7965 8134 8017 8186
rect 8029 8134 8081 8186
rect 8093 8134 8145 8186
rect 8157 8134 8209 8186
rect 8221 8134 8273 8186
rect 10771 8134 10823 8186
rect 10835 8134 10887 8186
rect 10899 8134 10951 8186
rect 10963 8134 11015 8186
rect 11027 8134 11079 8186
rect 1308 8032 1360 8084
rect 3056 8032 3108 8084
rect 4988 8032 5040 8084
rect 5448 8032 5500 8084
rect 6828 8075 6880 8084
rect 6828 8041 6837 8075
rect 6837 8041 6871 8075
rect 6871 8041 6880 8075
rect 6828 8032 6880 8041
rect 10416 8075 10468 8084
rect 10416 8041 10425 8075
rect 10425 8041 10459 8075
rect 10459 8041 10468 8075
rect 10416 8032 10468 8041
rect 2964 7964 3016 8016
rect 4068 7964 4120 8016
rect 7472 7964 7524 8016
rect 8208 8007 8260 8016
rect 8208 7973 8217 8007
rect 8217 7973 8251 8007
rect 8251 7973 8260 8007
rect 8208 7964 8260 7973
rect 1584 7828 1636 7880
rect 4528 7896 4580 7948
rect 6184 7896 6236 7948
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4252 7871 4304 7880
rect 4252 7837 4261 7871
rect 4261 7837 4295 7871
rect 4295 7837 4304 7871
rect 4252 7828 4304 7837
rect 6552 7828 6604 7880
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 7104 7760 7156 7812
rect 9128 7760 9180 7812
rect 2780 7692 2832 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 6828 7692 6880 7744
rect 3013 7590 3065 7642
rect 3077 7590 3129 7642
rect 3141 7590 3193 7642
rect 3205 7590 3257 7642
rect 3269 7590 3321 7642
rect 5819 7590 5871 7642
rect 5883 7590 5935 7642
rect 5947 7590 5999 7642
rect 6011 7590 6063 7642
rect 6075 7590 6127 7642
rect 8625 7590 8677 7642
rect 8689 7590 8741 7642
rect 8753 7590 8805 7642
rect 8817 7590 8869 7642
rect 8881 7590 8933 7642
rect 11431 7590 11483 7642
rect 11495 7590 11547 7642
rect 11559 7590 11611 7642
rect 11623 7590 11675 7642
rect 11687 7590 11739 7642
rect 4068 7420 4120 7472
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 3976 7259 4028 7268
rect 3976 7225 3985 7259
rect 3985 7225 4019 7259
rect 4019 7225 4028 7259
rect 3976 7216 4028 7225
rect 2688 7148 2740 7200
rect 4896 7352 4948 7404
rect 5540 7352 5592 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 6920 7488 6972 7540
rect 8208 7488 8260 7540
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 6736 7284 6788 7336
rect 8208 7352 8260 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 8668 7488 8720 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 10048 7488 10100 7540
rect 10508 7488 10560 7540
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 9588 7395 9640 7404
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 9588 7352 9640 7361
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 9772 7284 9824 7336
rect 10416 7284 10468 7336
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 10784 7395 10836 7404
rect 10784 7361 10793 7395
rect 10793 7361 10827 7395
rect 10827 7361 10836 7395
rect 10784 7352 10836 7361
rect 7104 7148 7156 7200
rect 7840 7148 7892 7200
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 2353 7046 2405 7098
rect 2417 7046 2469 7098
rect 2481 7046 2533 7098
rect 2545 7046 2597 7098
rect 2609 7046 2661 7098
rect 5159 7046 5211 7098
rect 5223 7046 5275 7098
rect 5287 7046 5339 7098
rect 5351 7046 5403 7098
rect 5415 7046 5467 7098
rect 7965 7046 8017 7098
rect 8029 7046 8081 7098
rect 8093 7046 8145 7098
rect 8157 7046 8209 7098
rect 8221 7046 8273 7098
rect 10771 7046 10823 7098
rect 10835 7046 10887 7098
rect 10899 7046 10951 7098
rect 10963 7046 11015 7098
rect 11027 7046 11079 7098
rect 6552 6944 6604 6996
rect 8392 6944 8444 6996
rect 2688 6808 2740 6860
rect 4528 6851 4580 6860
rect 4528 6817 4537 6851
rect 4537 6817 4571 6851
rect 4571 6817 4580 6851
rect 4528 6808 4580 6817
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 3792 6740 3844 6792
rect 3976 6740 4028 6792
rect 6184 6876 6236 6928
rect 8760 6876 8812 6928
rect 6644 6808 6696 6860
rect 9680 6944 9732 6996
rect 9772 6987 9824 6996
rect 9772 6953 9781 6987
rect 9781 6953 9815 6987
rect 9815 6953 9824 6987
rect 9772 6944 9824 6953
rect 10324 6987 10376 6996
rect 10324 6953 10333 6987
rect 10333 6953 10367 6987
rect 10367 6953 10376 6987
rect 10324 6944 10376 6953
rect 10692 6944 10744 6996
rect 9956 6876 10008 6928
rect 10416 6876 10468 6928
rect 9772 6808 9824 6860
rect 10876 6876 10928 6928
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 2872 6672 2924 6724
rect 6368 6672 6420 6724
rect 7196 6672 7248 6724
rect 7564 6672 7616 6724
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 8760 6740 8812 6792
rect 9680 6740 9732 6792
rect 10140 6740 10192 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 9772 6715 9824 6724
rect 9772 6681 9781 6715
rect 9781 6681 9815 6715
rect 9815 6681 9824 6715
rect 9772 6672 9824 6681
rect 2044 6604 2096 6656
rect 4068 6604 4120 6656
rect 4712 6647 4764 6656
rect 4712 6613 4721 6647
rect 4721 6613 4755 6647
rect 4755 6613 4764 6647
rect 4712 6604 4764 6613
rect 7288 6604 7340 6656
rect 9956 6647 10008 6656
rect 9956 6613 9965 6647
rect 9965 6613 9999 6647
rect 9999 6613 10008 6647
rect 9956 6604 10008 6613
rect 11244 6672 11296 6724
rect 11152 6604 11204 6656
rect 3013 6502 3065 6554
rect 3077 6502 3129 6554
rect 3141 6502 3193 6554
rect 3205 6502 3257 6554
rect 3269 6502 3321 6554
rect 5819 6502 5871 6554
rect 5883 6502 5935 6554
rect 5947 6502 5999 6554
rect 6011 6502 6063 6554
rect 6075 6502 6127 6554
rect 8625 6502 8677 6554
rect 8689 6502 8741 6554
rect 8753 6502 8805 6554
rect 8817 6502 8869 6554
rect 8881 6502 8933 6554
rect 11431 6502 11483 6554
rect 11495 6502 11547 6554
rect 11559 6502 11611 6554
rect 11623 6502 11675 6554
rect 11687 6502 11739 6554
rect 3976 6400 4028 6452
rect 8300 6400 8352 6452
rect 10692 6400 10744 6452
rect 11152 6400 11204 6452
rect 11244 6443 11296 6452
rect 11244 6409 11253 6443
rect 11253 6409 11287 6443
rect 11287 6409 11296 6443
rect 11244 6400 11296 6409
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 4068 6264 4120 6316
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 10048 6264 10100 6316
rect 1400 6128 1452 6180
rect 2872 6196 2924 6248
rect 4160 6196 4212 6248
rect 10692 6264 10744 6316
rect 10876 6264 10928 6316
rect 11336 6307 11388 6316
rect 11336 6273 11345 6307
rect 11345 6273 11379 6307
rect 11379 6273 11388 6307
rect 11336 6264 11388 6273
rect 1676 6060 1728 6112
rect 11888 6171 11940 6180
rect 11888 6137 11897 6171
rect 11897 6137 11931 6171
rect 11931 6137 11940 6171
rect 11888 6128 11940 6137
rect 2353 5958 2405 6010
rect 2417 5958 2469 6010
rect 2481 5958 2533 6010
rect 2545 5958 2597 6010
rect 2609 5958 2661 6010
rect 5159 5958 5211 6010
rect 5223 5958 5275 6010
rect 5287 5958 5339 6010
rect 5351 5958 5403 6010
rect 5415 5958 5467 6010
rect 7965 5958 8017 6010
rect 8029 5958 8081 6010
rect 8093 5958 8145 6010
rect 8157 5958 8209 6010
rect 8221 5958 8273 6010
rect 10771 5958 10823 6010
rect 10835 5958 10887 6010
rect 10899 5958 10951 6010
rect 10963 5958 11015 6010
rect 11027 5958 11079 6010
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 2964 5856 3016 5908
rect 8392 5856 8444 5908
rect 8668 5856 8720 5908
rect 10692 5899 10744 5908
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 4160 5720 4212 5772
rect 10048 5788 10100 5840
rect 11336 5788 11388 5840
rect 7288 5763 7340 5772
rect 7288 5729 7297 5763
rect 7297 5729 7331 5763
rect 7331 5729 7340 5763
rect 7288 5720 7340 5729
rect 1676 5695 1728 5704
rect 1676 5661 1710 5695
rect 1710 5661 1728 5695
rect 1676 5652 1728 5661
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 5632 5652 5684 5704
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 10508 5652 10560 5704
rect 10692 5652 10744 5704
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 4528 5584 4580 5636
rect 6184 5584 6236 5636
rect 6368 5627 6420 5636
rect 6368 5593 6377 5627
rect 6377 5593 6411 5627
rect 6411 5593 6420 5627
rect 6368 5584 6420 5593
rect 8300 5584 8352 5636
rect 5632 5559 5684 5568
rect 5632 5525 5641 5559
rect 5641 5525 5675 5559
rect 5675 5525 5684 5559
rect 5632 5516 5684 5525
rect 3013 5414 3065 5466
rect 3077 5414 3129 5466
rect 3141 5414 3193 5466
rect 3205 5414 3257 5466
rect 3269 5414 3321 5466
rect 5819 5414 5871 5466
rect 5883 5414 5935 5466
rect 5947 5414 5999 5466
rect 6011 5414 6063 5466
rect 6075 5414 6127 5466
rect 8625 5414 8677 5466
rect 8689 5414 8741 5466
rect 8753 5414 8805 5466
rect 8817 5414 8869 5466
rect 8881 5414 8933 5466
rect 11431 5414 11483 5466
rect 11495 5414 11547 5466
rect 11559 5414 11611 5466
rect 11623 5414 11675 5466
rect 11687 5414 11739 5466
rect 4068 5312 4120 5364
rect 4620 5244 4672 5296
rect 5724 5312 5776 5364
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 8300 5312 8352 5364
rect 7748 5244 7800 5296
rect 3976 5151 4028 5160
rect 3976 5117 3985 5151
rect 3985 5117 4019 5151
rect 4019 5117 4028 5151
rect 3976 5108 4028 5117
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 6920 5176 6972 5228
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 5724 5108 5776 5117
rect 7380 5108 7432 5160
rect 10508 5108 10560 5160
rect 4160 4972 4212 5024
rect 10692 4972 10744 5024
rect 2353 4870 2405 4922
rect 2417 4870 2469 4922
rect 2481 4870 2533 4922
rect 2545 4870 2597 4922
rect 2609 4870 2661 4922
rect 5159 4870 5211 4922
rect 5223 4870 5275 4922
rect 5287 4870 5339 4922
rect 5351 4870 5403 4922
rect 5415 4870 5467 4922
rect 7965 4870 8017 4922
rect 8029 4870 8081 4922
rect 8093 4870 8145 4922
rect 8157 4870 8209 4922
rect 8221 4870 8273 4922
rect 10771 4870 10823 4922
rect 10835 4870 10887 4922
rect 10899 4870 10951 4922
rect 10963 4870 11015 4922
rect 11027 4870 11079 4922
rect 3976 4768 4028 4820
rect 4620 4743 4672 4752
rect 4620 4709 4629 4743
rect 4629 4709 4663 4743
rect 4663 4709 4672 4743
rect 4620 4700 4672 4709
rect 4068 4564 4120 4616
rect 4712 4564 4764 4616
rect 5540 4768 5592 4820
rect 9036 4768 9088 4820
rect 9588 4768 9640 4820
rect 8392 4700 8444 4752
rect 10692 4700 10744 4752
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 5632 4564 5684 4616
rect 9036 4564 9088 4616
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 10692 4564 10744 4616
rect 3884 4496 3936 4548
rect 5724 4496 5776 4548
rect 6920 4496 6972 4548
rect 7564 4496 7616 4548
rect 10140 4496 10192 4548
rect 6184 4428 6236 4480
rect 8300 4428 8352 4480
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 9680 4428 9732 4480
rect 11244 4539 11296 4548
rect 11244 4505 11253 4539
rect 11253 4505 11287 4539
rect 11287 4505 11296 4539
rect 11244 4496 11296 4505
rect 3013 4326 3065 4378
rect 3077 4326 3129 4378
rect 3141 4326 3193 4378
rect 3205 4326 3257 4378
rect 3269 4326 3321 4378
rect 5819 4326 5871 4378
rect 5883 4326 5935 4378
rect 5947 4326 5999 4378
rect 6011 4326 6063 4378
rect 6075 4326 6127 4378
rect 8625 4326 8677 4378
rect 8689 4326 8741 4378
rect 8753 4326 8805 4378
rect 8817 4326 8869 4378
rect 8881 4326 8933 4378
rect 11431 4326 11483 4378
rect 11495 4326 11547 4378
rect 11559 4326 11611 4378
rect 11623 4326 11675 4378
rect 11687 4326 11739 4378
rect 4712 4224 4764 4276
rect 8392 4224 8444 4276
rect 9312 4224 9364 4276
rect 2136 4088 2188 4140
rect 2964 4088 3016 4140
rect 6184 4088 6236 4140
rect 2688 3952 2740 4004
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 6828 4156 6880 4208
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 9036 4156 9088 4208
rect 10232 4156 10284 4208
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8944 4088 8996 4140
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 7840 4020 7892 4072
rect 10416 4063 10468 4072
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10416 4020 10468 4029
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 11244 4088 11296 4140
rect 6092 3952 6144 4004
rect 7564 3952 7616 4004
rect 9956 3952 10008 4004
rect 10232 3952 10284 4004
rect 1768 3884 1820 3936
rect 6460 3884 6512 3936
rect 7472 3884 7524 3936
rect 10600 3884 10652 3936
rect 11612 3884 11664 3936
rect 2353 3782 2405 3834
rect 2417 3782 2469 3834
rect 2481 3782 2533 3834
rect 2545 3782 2597 3834
rect 2609 3782 2661 3834
rect 5159 3782 5211 3834
rect 5223 3782 5275 3834
rect 5287 3782 5339 3834
rect 5351 3782 5403 3834
rect 5415 3782 5467 3834
rect 7965 3782 8017 3834
rect 8029 3782 8081 3834
rect 8093 3782 8145 3834
rect 8157 3782 8209 3834
rect 8221 3782 8273 3834
rect 10771 3782 10823 3834
rect 10835 3782 10887 3834
rect 10899 3782 10951 3834
rect 10963 3782 11015 3834
rect 11027 3782 11079 3834
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 3884 3680 3936 3732
rect 1400 3544 1452 3596
rect 4160 3544 4212 3596
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 3608 3476 3660 3528
rect 5632 3476 5684 3528
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 6920 3680 6972 3732
rect 7656 3680 7708 3732
rect 7932 3680 7984 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 9680 3680 9732 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 2136 3451 2188 3460
rect 2136 3417 2145 3451
rect 2145 3417 2179 3451
rect 2179 3417 2188 3451
rect 2136 3408 2188 3417
rect 3700 3408 3752 3460
rect 6092 3408 6144 3460
rect 6828 3476 6880 3528
rect 7288 3544 7340 3596
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 1676 3340 1728 3392
rect 6276 3383 6328 3392
rect 6276 3349 6285 3383
rect 6285 3349 6319 3383
rect 6319 3349 6328 3383
rect 6276 3340 6328 3349
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 7748 3340 7800 3392
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 9772 3612 9824 3664
rect 10600 3612 10652 3664
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 11612 3476 11664 3528
rect 11888 3451 11940 3460
rect 11888 3417 11897 3451
rect 11897 3417 11931 3451
rect 11931 3417 11940 3451
rect 11888 3408 11940 3417
rect 3013 3238 3065 3290
rect 3077 3238 3129 3290
rect 3141 3238 3193 3290
rect 3205 3238 3257 3290
rect 3269 3238 3321 3290
rect 5819 3238 5871 3290
rect 5883 3238 5935 3290
rect 5947 3238 5999 3290
rect 6011 3238 6063 3290
rect 6075 3238 6127 3290
rect 8625 3238 8677 3290
rect 8689 3238 8741 3290
rect 8753 3238 8805 3290
rect 8817 3238 8869 3290
rect 8881 3238 8933 3290
rect 11431 3238 11483 3290
rect 11495 3238 11547 3290
rect 11559 3238 11611 3290
rect 11623 3238 11675 3290
rect 11687 3238 11739 3290
rect 2136 3136 2188 3188
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 6276 3136 6328 3188
rect 6920 3136 6972 3188
rect 7196 3136 7248 3188
rect 7932 3136 7984 3188
rect 9036 3136 9088 3188
rect 9404 3136 9456 3188
rect 7288 3111 7340 3120
rect 7288 3077 7297 3111
rect 7297 3077 7331 3111
rect 7331 3077 7340 3111
rect 7288 3068 7340 3077
rect 8024 3068 8076 3120
rect 9680 3068 9732 3120
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 1676 3043 1728 3052
rect 1676 3009 1710 3043
rect 1710 3009 1728 3043
rect 1676 3000 1728 3009
rect 4068 3000 4120 3052
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5540 3000 5592 3052
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10416 3000 10468 3052
rect 5632 2932 5684 2984
rect 6828 2932 6880 2984
rect 10600 2975 10652 2984
rect 10600 2941 10609 2975
rect 10609 2941 10643 2975
rect 10643 2941 10652 2975
rect 10600 2932 10652 2941
rect 6184 2796 6236 2848
rect 9680 2796 9732 2848
rect 2353 2694 2405 2746
rect 2417 2694 2469 2746
rect 2481 2694 2533 2746
rect 2545 2694 2597 2746
rect 2609 2694 2661 2746
rect 5159 2694 5211 2746
rect 5223 2694 5275 2746
rect 5287 2694 5339 2746
rect 5351 2694 5403 2746
rect 5415 2694 5467 2746
rect 7965 2694 8017 2746
rect 8029 2694 8081 2746
rect 8093 2694 8145 2746
rect 8157 2694 8209 2746
rect 8221 2694 8273 2746
rect 10771 2694 10823 2746
rect 10835 2694 10887 2746
rect 10899 2694 10951 2746
rect 10963 2694 11015 2746
rect 11027 2694 11079 2746
rect 5540 2592 5592 2644
rect 6184 2592 6236 2644
rect 7380 2456 7432 2508
rect 4068 2388 4120 2440
rect 5724 2388 5776 2440
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 7656 2388 7708 2440
rect 6460 2252 6512 2304
rect 7104 2252 7156 2304
rect 7748 2252 7800 2304
rect 3013 2150 3065 2202
rect 3077 2150 3129 2202
rect 3141 2150 3193 2202
rect 3205 2150 3257 2202
rect 3269 2150 3321 2202
rect 5819 2150 5871 2202
rect 5883 2150 5935 2202
rect 5947 2150 5999 2202
rect 6011 2150 6063 2202
rect 6075 2150 6127 2202
rect 8625 2150 8677 2202
rect 8689 2150 8741 2202
rect 8753 2150 8805 2202
rect 8817 2150 8869 2202
rect 8881 2150 8933 2202
rect 11431 2150 11483 2202
rect 11495 2150 11547 2202
rect 11559 2150 11611 2202
rect 11623 2150 11675 2202
rect 11687 2150 11739 2202
<< metal2 >>
rect 5814 14843 5870 15643
rect 6458 14843 6514 15643
rect 7102 14843 7158 15643
rect 7746 14843 7802 15643
rect 8390 14843 8446 15643
rect 5828 13274 5856 14843
rect 5736 13246 5856 13274
rect 3013 13084 3321 13093
rect 3013 13082 3019 13084
rect 3075 13082 3099 13084
rect 3155 13082 3179 13084
rect 3235 13082 3259 13084
rect 3315 13082 3321 13084
rect 3075 13030 3077 13082
rect 3257 13030 3259 13082
rect 3013 13028 3019 13030
rect 3075 13028 3099 13030
rect 3155 13028 3179 13030
rect 3235 13028 3259 13030
rect 3315 13028 3321 13030
rect 3013 13019 3321 13028
rect 5736 12986 5764 13246
rect 5819 13084 6127 13093
rect 5819 13082 5825 13084
rect 5881 13082 5905 13084
rect 5961 13082 5985 13084
rect 6041 13082 6065 13084
rect 6121 13082 6127 13084
rect 5881 13030 5883 13082
rect 6063 13030 6065 13082
rect 5819 13028 5825 13030
rect 5881 13028 5905 13030
rect 5961 13028 5985 13030
rect 6041 13028 6065 13030
rect 6121 13028 6127 13030
rect 5819 13019 6127 13028
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 6472 12918 6500 14843
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 7116 12850 7144 14843
rect 7760 12850 7788 14843
rect 8404 12850 8432 14843
rect 8625 13084 8933 13093
rect 8625 13082 8631 13084
rect 8687 13082 8711 13084
rect 8767 13082 8791 13084
rect 8847 13082 8871 13084
rect 8927 13082 8933 13084
rect 8687 13030 8689 13082
rect 8869 13030 8871 13082
rect 8625 13028 8631 13030
rect 8687 13028 8711 13030
rect 8767 13028 8791 13030
rect 8847 13028 8871 13030
rect 8927 13028 8933 13030
rect 8625 13019 8933 13028
rect 11431 13084 11739 13093
rect 11431 13082 11437 13084
rect 11493 13082 11517 13084
rect 11573 13082 11597 13084
rect 11653 13082 11677 13084
rect 11733 13082 11739 13084
rect 11493 13030 11495 13082
rect 11675 13030 11677 13082
rect 11431 13028 11437 13030
rect 11493 13028 11517 13030
rect 11573 13028 11597 13030
rect 11653 13028 11677 13030
rect 11733 13028 11739 13030
rect 11431 13019 11739 13028
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 2353 12540 2661 12549
rect 2353 12538 2359 12540
rect 2415 12538 2439 12540
rect 2495 12538 2519 12540
rect 2575 12538 2599 12540
rect 2655 12538 2661 12540
rect 2415 12486 2417 12538
rect 2597 12486 2599 12538
rect 2353 12484 2359 12486
rect 2415 12484 2439 12486
rect 2495 12484 2519 12486
rect 2575 12484 2599 12486
rect 2655 12484 2661 12486
rect 2353 12475 2661 12484
rect 5159 12540 5467 12549
rect 5159 12538 5165 12540
rect 5221 12538 5245 12540
rect 5301 12538 5325 12540
rect 5381 12538 5405 12540
rect 5461 12538 5467 12540
rect 5221 12486 5223 12538
rect 5403 12486 5405 12538
rect 5159 12484 5165 12486
rect 5221 12484 5245 12486
rect 5301 12484 5325 12486
rect 5381 12484 5405 12486
rect 5461 12484 5467 12486
rect 5159 12475 5467 12484
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 1584 12164 1636 12170
rect 1584 12106 1636 12112
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1596 11082 1624 12106
rect 2332 11898 2360 12106
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2608 11762 2636 12242
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 3013 11996 3321 12005
rect 3013 11994 3019 11996
rect 3075 11994 3099 11996
rect 3155 11994 3179 11996
rect 3235 11994 3259 11996
rect 3315 11994 3321 11996
rect 3075 11942 3077 11994
rect 3257 11942 3259 11994
rect 3013 11940 3019 11942
rect 3075 11940 3099 11942
rect 3155 11940 3179 11942
rect 3235 11940 3259 11942
rect 3315 11940 3321 11942
rect 3013 11931 3321 11940
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2608 11642 2636 11698
rect 2608 11614 2728 11642
rect 2353 11452 2661 11461
rect 2353 11450 2359 11452
rect 2415 11450 2439 11452
rect 2495 11450 2519 11452
rect 2575 11450 2599 11452
rect 2655 11450 2661 11452
rect 2415 11398 2417 11450
rect 2597 11398 2599 11450
rect 2353 11396 2359 11398
rect 2415 11396 2439 11398
rect 2495 11396 2519 11398
rect 2575 11396 2599 11398
rect 2655 11396 2661 11398
rect 2353 11387 2661 11396
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1306 10296 1362 10305
rect 1306 10231 1308 10240
rect 1360 10231 1362 10240
rect 1308 10202 1360 10208
rect 1412 9518 1440 10542
rect 1596 10062 1624 11018
rect 2353 10364 2661 10373
rect 2353 10362 2359 10364
rect 2415 10362 2439 10364
rect 2495 10362 2519 10364
rect 2575 10362 2599 10364
rect 2655 10362 2661 10364
rect 2415 10310 2417 10362
rect 2597 10310 2599 10362
rect 2353 10308 2359 10310
rect 2415 10308 2439 10310
rect 2495 10308 2519 10310
rect 2575 10308 2599 10310
rect 2655 10308 2661 10310
rect 2353 10299 2661 10308
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 2700 9518 2728 11614
rect 2792 11286 2820 11766
rect 3344 11354 3372 11766
rect 4540 11354 4568 12106
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 4724 11150 4752 11494
rect 4908 11354 4936 11698
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5000 11218 5028 12174
rect 5552 12170 5580 12786
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5552 11898 5580 12106
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5540 11756 5592 11762
rect 5644 11744 5672 12038
rect 5819 11996 6127 12005
rect 5819 11994 5825 11996
rect 5881 11994 5905 11996
rect 5961 11994 5985 11996
rect 6041 11994 6065 11996
rect 6121 11994 6127 11996
rect 5881 11942 5883 11994
rect 6063 11942 6065 11994
rect 5819 11940 5825 11942
rect 5881 11940 5905 11942
rect 5961 11940 5985 11942
rect 6041 11940 6065 11942
rect 6121 11940 6127 11942
rect 5819 11931 6127 11940
rect 6196 11830 6224 12310
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 5592 11716 5672 11744
rect 5540 11698 5592 11704
rect 5159 11452 5467 11461
rect 5159 11450 5165 11452
rect 5221 11450 5245 11452
rect 5301 11450 5325 11452
rect 5381 11450 5405 11452
rect 5461 11450 5467 11452
rect 5221 11398 5223 11450
rect 5403 11398 5405 11450
rect 5159 11396 5165 11398
rect 5221 11396 5245 11398
rect 5301 11396 5325 11398
rect 5381 11396 5405 11398
rect 5461 11396 5467 11398
rect 5159 11387 5467 11396
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 3013 10908 3321 10917
rect 3013 10906 3019 10908
rect 3075 10906 3099 10908
rect 3155 10906 3179 10908
rect 3235 10906 3259 10908
rect 3315 10906 3321 10908
rect 3075 10854 3077 10906
rect 3257 10854 3259 10906
rect 3013 10852 3019 10854
rect 3075 10852 3099 10854
rect 3155 10852 3179 10854
rect 3235 10852 3259 10854
rect 3315 10852 3321 10854
rect 3013 10843 3321 10852
rect 3436 10674 3464 11086
rect 5000 11082 5028 11154
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3013 9820 3321 9829
rect 3013 9818 3019 9820
rect 3075 9818 3099 9820
rect 3155 9818 3179 9820
rect 3235 9818 3259 9820
rect 3315 9818 3321 9820
rect 3075 9766 3077 9818
rect 3257 9766 3259 9818
rect 3013 9764 3019 9766
rect 3075 9764 3099 9766
rect 3155 9764 3179 9766
rect 3235 9764 3259 9766
rect 3315 9764 3321 9766
rect 3013 9755 3321 9764
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 1688 9178 1716 9454
rect 2700 9382 2728 9454
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2353 9276 2661 9285
rect 2353 9274 2359 9276
rect 2415 9274 2439 9276
rect 2495 9274 2519 9276
rect 2575 9274 2599 9276
rect 2655 9274 2661 9276
rect 2415 9222 2417 9274
rect 2597 9222 2599 9274
rect 2353 9220 2359 9222
rect 2415 9220 2439 9222
rect 2495 9220 2519 9222
rect 2575 9220 2599 9222
rect 2655 9220 2661 9222
rect 2353 9211 2661 9220
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 2700 9042 2728 9318
rect 2792 9178 2820 9522
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2700 8634 2728 8978
rect 3436 8974 3464 10610
rect 5000 9738 5028 11018
rect 5092 10266 5120 11086
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 10810 5396 10950
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5644 10674 5672 11716
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5159 10364 5467 10373
rect 5159 10362 5165 10364
rect 5221 10362 5245 10364
rect 5301 10362 5325 10364
rect 5381 10362 5405 10364
rect 5461 10362 5467 10364
rect 5221 10310 5223 10362
rect 5403 10310 5405 10362
rect 5159 10308 5165 10310
rect 5221 10308 5245 10310
rect 5301 10308 5325 10310
rect 5381 10308 5405 10310
rect 5461 10308 5467 10310
rect 5159 10299 5467 10308
rect 5552 10266 5580 10542
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 4908 9710 5028 9738
rect 4908 8974 4936 9710
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 3013 8732 3321 8741
rect 3013 8730 3019 8732
rect 3075 8730 3099 8732
rect 3155 8730 3179 8732
rect 3235 8730 3259 8732
rect 3315 8730 3321 8732
rect 3075 8678 3077 8730
rect 3257 8678 3259 8730
rect 3013 8676 3019 8678
rect 3075 8676 3099 8678
rect 3155 8676 3179 8678
rect 3235 8676 3259 8678
rect 3315 8676 3321 8678
rect 3013 8667 3321 8676
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 1584 8288 1636 8294
rect 1306 8256 1362 8265
rect 1584 8230 1636 8236
rect 1306 8191 1362 8200
rect 1320 8090 1348 8191
rect 1308 8084 1360 8090
rect 1308 8026 1360 8032
rect 1596 7886 1624 8230
rect 2353 8188 2661 8197
rect 2353 8186 2359 8188
rect 2415 8186 2439 8188
rect 2495 8186 2519 8188
rect 2575 8186 2599 8188
rect 2655 8186 2661 8188
rect 2415 8134 2417 8186
rect 2597 8134 2599 8186
rect 2353 8132 2359 8134
rect 2415 8132 2439 8134
rect 2495 8132 2519 8134
rect 2575 8132 2599 8134
rect 2655 8132 2661 8134
rect 2353 8123 2661 8132
rect 2976 8022 3004 8366
rect 3068 8090 3096 8366
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 3804 7886 3832 8910
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4250 8256 4306 8265
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2353 7100 2661 7109
rect 2353 7098 2359 7100
rect 2415 7098 2439 7100
rect 2495 7098 2519 7100
rect 2575 7098 2599 7100
rect 2655 7098 2661 7100
rect 2415 7046 2417 7098
rect 2597 7046 2599 7098
rect 2353 7044 2359 7046
rect 2415 7044 2439 7046
rect 2495 7044 2519 7046
rect 2575 7044 2599 7046
rect 2655 7044 2661 7046
rect 2353 7035 2661 7044
rect 2700 6866 2728 7142
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 6322 2084 6598
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1400 6180 1452 6186
rect 1400 6122 1452 6128
rect 1412 5778 1440 6122
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1688 5710 1716 6054
rect 2353 6012 2661 6021
rect 2353 6010 2359 6012
rect 2415 6010 2439 6012
rect 2495 6010 2519 6012
rect 2575 6010 2599 6012
rect 2655 6010 2661 6012
rect 2415 5958 2417 6010
rect 2597 5958 2599 6010
rect 2353 5956 2359 5958
rect 2415 5956 2439 5958
rect 2495 5956 2519 5958
rect 2575 5956 2599 5958
rect 2655 5956 2661 5958
rect 2353 5947 2661 5956
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 2353 4924 2661 4933
rect 2353 4922 2359 4924
rect 2415 4922 2439 4924
rect 2495 4922 2519 4924
rect 2575 4922 2599 4924
rect 2655 4922 2661 4924
rect 2415 4870 2417 4922
rect 2597 4870 2599 4922
rect 2353 4868 2359 4870
rect 2415 4868 2439 4870
rect 2495 4868 2519 4870
rect 2575 4868 2599 4870
rect 2655 4868 2661 4870
rect 2353 4859 2661 4868
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 3058 1440 3538
rect 1780 3534 1808 3878
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2148 3466 2176 4082
rect 2700 4010 2728 6802
rect 2792 6798 2820 7686
rect 3013 7644 3321 7653
rect 3013 7642 3019 7644
rect 3075 7642 3099 7644
rect 3155 7642 3179 7644
rect 3235 7642 3259 7644
rect 3315 7642 3321 7644
rect 3075 7590 3077 7642
rect 3257 7590 3259 7642
rect 3013 7588 3019 7590
rect 3075 7588 3099 7590
rect 3155 7588 3179 7590
rect 3235 7588 3259 7590
rect 3315 7588 3321 7590
rect 3013 7579 3321 7588
rect 3804 6798 3832 7822
rect 4080 7478 4108 7958
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 2792 5794 2820 6734
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2884 6254 2912 6666
rect 3013 6556 3321 6565
rect 3013 6554 3019 6556
rect 3075 6554 3099 6556
rect 3155 6554 3179 6556
rect 3235 6554 3259 6556
rect 3315 6554 3321 6556
rect 3075 6502 3077 6554
rect 3257 6502 3259 6554
rect 3013 6500 3019 6502
rect 3075 6500 3099 6502
rect 3155 6500 3179 6502
rect 3235 6500 3259 6502
rect 3315 6500 3321 6502
rect 3013 6491 3321 6500
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2884 5914 2912 6190
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2976 5794 3004 5850
rect 2792 5766 3004 5794
rect 2792 4162 2820 5766
rect 3013 5468 3321 5477
rect 3013 5466 3019 5468
rect 3075 5466 3099 5468
rect 3155 5466 3179 5468
rect 3235 5466 3259 5468
rect 3315 5466 3321 5468
rect 3075 5414 3077 5466
rect 3257 5414 3259 5466
rect 3013 5412 3019 5414
rect 3075 5412 3099 5414
rect 3155 5412 3179 5414
rect 3235 5412 3259 5414
rect 3315 5412 3321 5414
rect 3013 5403 3321 5412
rect 3896 4554 3924 7346
rect 4068 7336 4120 7342
rect 4172 7290 4200 8230
rect 4250 8191 4306 8200
rect 4264 7886 4292 8191
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4120 7284 4200 7290
rect 4068 7278 4200 7284
rect 3976 7268 4028 7274
rect 4080 7262 4200 7278
rect 3976 7210 4028 7216
rect 3988 6798 4016 7210
rect 4540 6866 4568 7890
rect 4908 7410 4936 8910
rect 5000 8090 5028 9522
rect 5092 8294 5120 9930
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5159 9276 5467 9285
rect 5159 9274 5165 9276
rect 5221 9274 5245 9276
rect 5301 9274 5325 9276
rect 5381 9274 5405 9276
rect 5461 9274 5467 9276
rect 5221 9222 5223 9274
rect 5403 9222 5405 9274
rect 5159 9220 5165 9222
rect 5221 9220 5245 9222
rect 5301 9220 5325 9222
rect 5381 9220 5405 9222
rect 5461 9220 5467 9222
rect 5159 9211 5467 9220
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 8498 5304 8910
rect 5552 8906 5580 9318
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5552 8498 5580 8842
rect 5644 8498 5672 10610
rect 5736 10538 5764 11086
rect 5819 10908 6127 10917
rect 5819 10906 5825 10908
rect 5881 10906 5905 10908
rect 5961 10906 5985 10908
rect 6041 10906 6065 10908
rect 6121 10906 6127 10908
rect 5881 10854 5883 10906
rect 6063 10854 6065 10906
rect 5819 10852 5825 10854
rect 5881 10852 5905 10854
rect 5961 10852 5985 10854
rect 6041 10852 6065 10854
rect 6121 10852 6127 10854
rect 5819 10843 6127 10852
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5920 10418 5948 10474
rect 5920 10390 6040 10418
rect 6012 10198 6040 10390
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 6012 10062 6040 10134
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5819 9820 6127 9829
rect 5819 9818 5825 9820
rect 5881 9818 5905 9820
rect 5961 9818 5985 9820
rect 6041 9818 6065 9820
rect 6121 9818 6127 9820
rect 5881 9766 5883 9818
rect 6063 9766 6065 9818
rect 5819 9764 5825 9766
rect 5881 9764 5905 9766
rect 5961 9764 5985 9766
rect 6041 9764 6065 9766
rect 6121 9764 6127 9766
rect 5819 9755 6127 9764
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9178 5948 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5736 8634 5764 8978
rect 5819 8732 6127 8741
rect 5819 8730 5825 8732
rect 5881 8730 5905 8732
rect 5961 8730 5985 8732
rect 6041 8730 6065 8732
rect 6121 8730 6127 8732
rect 5881 8678 5883 8730
rect 6063 8678 6065 8730
rect 5819 8676 5825 8678
rect 5881 8676 5905 8678
rect 5961 8676 5985 8678
rect 6041 8676 6065 8678
rect 6121 8676 6127 8678
rect 5819 8667 6127 8676
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5159 8188 5467 8197
rect 5159 8186 5165 8188
rect 5221 8186 5245 8188
rect 5301 8186 5325 8188
rect 5381 8186 5405 8188
rect 5461 8186 5467 8188
rect 5221 8134 5223 8186
rect 5403 8134 5405 8186
rect 5159 8132 5165 8134
rect 5221 8132 5245 8134
rect 5301 8132 5325 8134
rect 5381 8132 5405 8134
rect 5461 8132 5467 8134
rect 5159 8123 5467 8132
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 5460 7188 5488 8026
rect 5552 7410 5580 8298
rect 6196 7954 6224 11562
rect 6380 10810 6408 11698
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6656 11150 6684 11562
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6564 10674 6592 11086
rect 6932 10742 6960 12786
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11898 7420 12174
rect 7576 12170 7604 12582
rect 7965 12540 8273 12549
rect 7965 12538 7971 12540
rect 8027 12538 8051 12540
rect 8107 12538 8131 12540
rect 8187 12538 8211 12540
rect 8267 12538 8273 12540
rect 8027 12486 8029 12538
rect 8209 12486 8211 12538
rect 7965 12484 7971 12486
rect 8027 12484 8051 12486
rect 8107 12484 8131 12486
rect 8187 12484 8211 12486
rect 8267 12484 8273 12486
rect 7965 12475 8273 12484
rect 8312 12238 8340 12582
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 8634 6408 9930
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9586 6500 9862
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6472 7698 6500 9522
rect 6564 9518 6592 10610
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 9586 6868 10542
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 7024 8838 7052 11290
rect 7300 9654 7328 11630
rect 7392 11082 7420 11630
rect 7484 11354 7512 11630
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7576 10674 7604 12106
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7760 11762 7788 12038
rect 7944 11830 7972 12038
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7760 11234 7788 11698
rect 8128 11694 8156 12038
rect 8312 11762 8340 12174
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 8404 11762 8432 12106
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8116 11688 8168 11694
rect 7668 11218 7788 11234
rect 7656 11212 7788 11218
rect 7708 11206 7788 11212
rect 7852 11636 8116 11642
rect 7852 11630 8168 11636
rect 7852 11614 8156 11630
rect 7656 11154 7708 11160
rect 7852 11150 7880 11614
rect 7965 11452 8273 11461
rect 7965 11450 7971 11452
rect 8027 11450 8051 11452
rect 8107 11450 8131 11452
rect 8187 11450 8211 11452
rect 8267 11450 8273 11452
rect 8027 11398 8029 11450
rect 8209 11398 8211 11450
rect 7965 11396 7971 11398
rect 8027 11396 8051 11398
rect 8107 11396 8131 11398
rect 8187 11396 8211 11398
rect 8267 11396 8273 11398
rect 7965 11387 8273 11396
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 8312 10470 8340 11698
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 11354 8432 11562
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 7965 10364 8273 10373
rect 7965 10362 7971 10364
rect 8027 10362 8051 10364
rect 8107 10362 8131 10364
rect 8187 10362 8211 10364
rect 8267 10362 8273 10364
rect 8027 10310 8029 10362
rect 8209 10310 8211 10362
rect 7965 10308 7971 10310
rect 8027 10308 8051 10310
rect 8107 10308 8131 10310
rect 8187 10308 8211 10310
rect 8267 10308 8273 10310
rect 7965 10299 8273 10308
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 9042 7512 9454
rect 7965 9276 8273 9285
rect 7965 9274 7971 9276
rect 8027 9274 8051 9276
rect 8107 9274 8131 9276
rect 8187 9274 8211 9276
rect 8267 9274 8273 9276
rect 8027 9222 8029 9274
rect 8209 9222 8211 9274
rect 7965 9220 7971 9222
rect 8027 9220 8051 9222
rect 8107 9220 8131 9222
rect 8187 9220 8211 9222
rect 8267 9220 8273 9222
rect 7965 9211 8273 9220
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7484 8906 7512 8978
rect 8312 8906 8340 9114
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6656 8294 6684 8502
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6564 7886 6592 8230
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6552 7744 6604 7750
rect 6472 7692 6552 7698
rect 6472 7686 6604 7692
rect 6472 7670 6592 7686
rect 5819 7644 6127 7653
rect 5819 7642 5825 7644
rect 5881 7642 5905 7644
rect 5961 7642 5985 7644
rect 6041 7642 6065 7644
rect 6121 7642 6127 7644
rect 5881 7590 5883 7642
rect 6063 7590 6065 7642
rect 5819 7588 5825 7590
rect 5881 7588 5905 7590
rect 5961 7588 5985 7590
rect 6041 7588 6065 7590
rect 6121 7588 6127 7590
rect 5819 7579 6127 7588
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 5460 7160 5580 7188
rect 5159 7100 5467 7109
rect 5159 7098 5165 7100
rect 5221 7098 5245 7100
rect 5301 7098 5325 7100
rect 5381 7098 5405 7100
rect 5461 7098 5467 7100
rect 5221 7046 5223 7098
rect 5403 7046 5405 7098
rect 5159 7044 5165 7046
rect 5221 7044 5245 7046
rect 5301 7044 5325 7046
rect 5381 7044 5405 7046
rect 5461 7044 5467 7046
rect 5159 7035 5467 7044
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 6458 4016 6734
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 4080 6322 4108 6598
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4080 5370 4108 6258
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4172 5778 4200 6190
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3988 4826 4016 5102
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4080 4622 4108 5306
rect 4172 5030 4200 5714
rect 4540 5642 4568 6802
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 3013 4380 3321 4389
rect 3013 4378 3019 4380
rect 3075 4378 3099 4380
rect 3155 4378 3179 4380
rect 3235 4378 3259 4380
rect 3315 4378 3321 4380
rect 3075 4326 3077 4378
rect 3257 4326 3259 4378
rect 3013 4324 3019 4326
rect 3075 4324 3099 4326
rect 3155 4324 3179 4326
rect 3235 4324 3259 4326
rect 3315 4324 3321 4326
rect 3013 4315 3321 4324
rect 2792 4146 3004 4162
rect 2792 4140 3016 4146
rect 2792 4134 2964 4140
rect 2964 4082 3016 4088
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2353 3836 2661 3845
rect 2353 3834 2359 3836
rect 2415 3834 2439 3836
rect 2495 3834 2519 3836
rect 2575 3834 2599 3836
rect 2655 3834 2661 3836
rect 2415 3782 2417 3834
rect 2597 3782 2599 3834
rect 2353 3780 2359 3782
rect 2415 3780 2439 3782
rect 2495 3780 2519 3782
rect 2575 3780 2599 3782
rect 2655 3780 2661 3782
rect 2353 3771 2661 3780
rect 3620 3738 3648 4014
rect 3896 3738 3924 4490
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3620 3534 3648 3674
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1688 3058 1716 3334
rect 2148 3194 2176 3402
rect 3013 3292 3321 3301
rect 3013 3290 3019 3292
rect 3075 3290 3099 3292
rect 3155 3290 3179 3292
rect 3235 3290 3259 3292
rect 3315 3290 3321 3292
rect 3075 3238 3077 3290
rect 3257 3238 3259 3290
rect 3013 3236 3019 3238
rect 3075 3236 3099 3238
rect 3155 3236 3179 3238
rect 3235 3236 3259 3238
rect 3315 3236 3321 3238
rect 3013 3227 3321 3236
rect 3712 3194 3740 3402
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 4080 3058 4108 4558
rect 4172 3602 4200 4966
rect 4632 4758 4660 5238
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4724 4622 4752 6598
rect 5159 6012 5467 6021
rect 5159 6010 5165 6012
rect 5221 6010 5245 6012
rect 5301 6010 5325 6012
rect 5381 6010 5405 6012
rect 5461 6010 5467 6012
rect 5221 5958 5223 6010
rect 5403 5958 5405 6010
rect 5159 5956 5165 5958
rect 5221 5956 5245 5958
rect 5301 5956 5325 5958
rect 5381 5956 5405 5958
rect 5461 5956 5467 5958
rect 5159 5947 5467 5956
rect 5552 5710 5580 7160
rect 5644 5710 5672 7346
rect 6196 6934 6224 7346
rect 6564 7002 6592 7346
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6656 6866 6684 8230
rect 6748 7342 6776 8434
rect 6840 8090 6868 8434
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6840 7410 6868 7686
rect 6932 7546 6960 7822
rect 7116 7818 7144 8434
rect 7484 8022 7512 8842
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6748 6798 6776 7278
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 5819 6556 6127 6565
rect 5819 6554 5825 6556
rect 5881 6554 5905 6556
rect 5961 6554 5985 6556
rect 6041 6554 6065 6556
rect 6121 6554 6127 6556
rect 5881 6502 5883 6554
rect 6063 6502 6065 6554
rect 5819 6500 5825 6502
rect 5881 6500 5905 6502
rect 5961 6500 5985 6502
rect 6041 6500 6065 6502
rect 6121 6500 6127 6502
rect 5819 6491 6127 6500
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5632 5704 5684 5710
rect 5684 5652 5764 5658
rect 5632 5646 5764 5652
rect 5644 5630 5764 5646
rect 6380 5642 6408 6666
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5159 4924 5467 4933
rect 5159 4922 5165 4924
rect 5221 4922 5245 4924
rect 5301 4922 5325 4924
rect 5381 4922 5405 4924
rect 5461 4922 5467 4924
rect 5221 4870 5223 4922
rect 5403 4870 5405 4922
rect 5159 4868 5165 4870
rect 5221 4868 5245 4870
rect 5301 4868 5325 4870
rect 5381 4868 5405 4870
rect 5461 4868 5467 4870
rect 5159 4859 5467 4868
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4282 4752 4558
rect 5552 4434 5580 4762
rect 5644 4622 5672 5510
rect 5736 5370 5764 5630
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 5819 5468 6127 5477
rect 5819 5466 5825 5468
rect 5881 5466 5905 5468
rect 5961 5466 5985 5468
rect 6041 5466 6065 5468
rect 6121 5466 6127 5468
rect 5881 5414 5883 5466
rect 6063 5414 6065 5466
rect 5819 5412 5825 5414
rect 5881 5412 5905 5414
rect 5961 5412 5985 5414
rect 6041 5412 6065 5414
rect 6121 5412 6127 5414
rect 5819 5403 6127 5412
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5736 4554 5764 5102
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 6196 4486 6224 5578
rect 6380 5370 6408 5578
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6184 4480 6236 4486
rect 5552 4406 5764 4434
rect 6184 4422 6236 4428
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 5159 3836 5467 3845
rect 5159 3834 5165 3836
rect 5221 3834 5245 3836
rect 5301 3834 5325 3836
rect 5381 3834 5405 3836
rect 5461 3834 5467 3836
rect 5221 3782 5223 3834
rect 5403 3782 5405 3834
rect 5159 3780 5165 3782
rect 5221 3780 5245 3782
rect 5301 3780 5325 3782
rect 5381 3780 5405 3782
rect 5461 3780 5467 3782
rect 5159 3771 5467 3780
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 3058 4200 3538
rect 5736 3534 5764 4406
rect 5819 4380 6127 4389
rect 5819 4378 5825 4380
rect 5881 4378 5905 4380
rect 5961 4378 5985 4380
rect 6041 4378 6065 4380
rect 6121 4378 6127 4380
rect 5881 4326 5883 4378
rect 6063 4326 6065 4378
rect 5819 4324 5825 4326
rect 5881 4324 5905 4326
rect 5961 4324 5985 4326
rect 6041 4324 6065 4326
rect 6121 4324 6127 4326
rect 5819 4315 6127 4324
rect 6196 4146 6224 4422
rect 6840 4214 6868 7346
rect 7116 7206 7144 7754
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7576 6730 7604 8774
rect 8220 8634 8248 8774
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 8430 8340 8842
rect 8404 8498 8432 11018
rect 8496 10742 8524 12582
rect 10771 12540 11079 12549
rect 10771 12538 10777 12540
rect 10833 12538 10857 12540
rect 10913 12538 10937 12540
rect 10993 12538 11017 12540
rect 11073 12538 11079 12540
rect 10833 12486 10835 12538
rect 11015 12486 11017 12538
rect 10771 12484 10777 12486
rect 10833 12484 10857 12486
rect 10913 12484 10937 12486
rect 10993 12484 11017 12486
rect 11073 12484 11079 12486
rect 10771 12475 11079 12484
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 8625 11996 8933 12005
rect 8625 11994 8631 11996
rect 8687 11994 8711 11996
rect 8767 11994 8791 11996
rect 8847 11994 8871 11996
rect 8927 11994 8933 11996
rect 8687 11942 8689 11994
rect 8869 11942 8871 11994
rect 8625 11940 8631 11942
rect 8687 11940 8711 11942
rect 8767 11940 8791 11942
rect 8847 11940 8871 11942
rect 8927 11940 8933 11942
rect 8625 11931 8933 11940
rect 9324 11898 9352 12038
rect 9876 11898 9904 12106
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10336 11762 10364 12174
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 8625 10908 8933 10917
rect 8625 10906 8631 10908
rect 8687 10906 8711 10908
rect 8767 10906 8791 10908
rect 8847 10906 8871 10908
rect 8927 10906 8933 10908
rect 8687 10854 8689 10906
rect 8869 10854 8871 10906
rect 8625 10852 8631 10854
rect 8687 10852 8711 10854
rect 8767 10852 8791 10854
rect 8847 10852 8871 10854
rect 8927 10852 8933 10854
rect 8625 10843 8933 10852
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8496 10062 8524 10678
rect 9876 10674 9904 11630
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8588 9994 8616 10610
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8625 9820 8933 9829
rect 8625 9818 8631 9820
rect 8687 9818 8711 9820
rect 8767 9818 8791 9820
rect 8847 9818 8871 9820
rect 8927 9818 8933 9820
rect 8687 9766 8689 9818
rect 8869 9766 8871 9818
rect 8625 9764 8631 9766
rect 8687 9764 8711 9766
rect 8767 9764 8791 9766
rect 8847 9764 8871 9766
rect 8927 9764 8933 9766
rect 8625 9755 8933 9764
rect 9140 9518 9168 10134
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9654 9352 9862
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9416 9586 9444 9930
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9140 9178 9168 9454
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9416 9042 9444 9522
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 8625 8732 8933 8741
rect 8625 8730 8631 8732
rect 8687 8730 8711 8732
rect 8767 8730 8791 8732
rect 8847 8730 8871 8732
rect 8927 8730 8933 8732
rect 8687 8678 8689 8730
rect 8869 8678 8871 8730
rect 8625 8676 8631 8678
rect 8687 8676 8711 8678
rect 8767 8676 8791 8678
rect 8847 8676 8871 8678
rect 8927 8676 8933 8678
rect 8625 8667 8933 8676
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 7965 8188 8273 8197
rect 7965 8186 7971 8188
rect 8027 8186 8051 8188
rect 8107 8186 8131 8188
rect 8187 8186 8211 8188
rect 8267 8186 8273 8188
rect 8027 8134 8029 8186
rect 8209 8134 8211 8186
rect 7965 8132 7971 8134
rect 8027 8132 8051 8134
rect 8107 8132 8131 8134
rect 8187 8132 8211 8134
rect 8267 8132 8273 8134
rect 7965 8123 8273 8132
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8220 7546 8248 7958
rect 8625 7644 8933 7653
rect 8625 7642 8631 7644
rect 8687 7642 8711 7644
rect 8767 7642 8791 7644
rect 8847 7642 8871 7644
rect 8927 7642 8933 7644
rect 8687 7590 8689 7642
rect 8869 7590 8871 7642
rect 8625 7588 8631 7590
rect 8687 7588 8711 7590
rect 8767 7588 8791 7590
rect 8847 7588 8871 7590
rect 8927 7588 8933 7590
rect 8625 7579 8933 7588
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8220 7290 8248 7346
rect 8220 7262 8340 7290
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 6798 7880 7142
rect 7965 7100 8273 7109
rect 7965 7098 7971 7100
rect 8027 7098 8051 7100
rect 8107 7098 8131 7100
rect 8187 7098 8211 7100
rect 8267 7098 8273 7100
rect 8027 7046 8029 7098
rect 8209 7046 8211 7098
rect 7965 7044 7971 7046
rect 8027 7044 8051 7046
rect 8107 7044 8131 7046
rect 8187 7044 8211 7046
rect 8267 7044 8273 7046
rect 7965 7035 8273 7044
rect 8312 6798 8340 7262
rect 8404 7002 8432 7346
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8680 6882 8708 7482
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8772 6934 8800 7346
rect 8404 6854 8708 6882
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6932 4554 6960 5170
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6932 4146 6960 4490
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 6104 3482 6132 3946
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3602 6500 3878
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6828 3528 6880 3534
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 2353 2748 2661 2757
rect 2353 2746 2359 2748
rect 2415 2746 2439 2748
rect 2495 2746 2519 2748
rect 2575 2746 2599 2748
rect 2655 2746 2661 2748
rect 2415 2694 2417 2746
rect 2597 2694 2599 2746
rect 2353 2692 2359 2694
rect 2415 2692 2439 2694
rect 2495 2692 2519 2694
rect 2575 2692 2599 2694
rect 2655 2692 2661 2694
rect 2353 2683 2661 2692
rect 4080 2446 4108 2994
rect 5159 2748 5467 2757
rect 5159 2746 5165 2748
rect 5221 2746 5245 2748
rect 5301 2746 5325 2748
rect 5381 2746 5405 2748
rect 5461 2746 5467 2748
rect 5221 2694 5223 2746
rect 5403 2694 5405 2746
rect 5159 2692 5165 2694
rect 5221 2692 5245 2694
rect 5301 2692 5325 2694
rect 5381 2692 5405 2694
rect 5461 2692 5467 2694
rect 5159 2683 5467 2692
rect 5552 2650 5580 2994
rect 5644 2990 5672 3470
rect 6104 3466 6224 3482
rect 6828 3470 6880 3476
rect 6092 3460 6224 3466
rect 6144 3454 6224 3460
rect 6092 3402 6144 3408
rect 5819 3292 6127 3301
rect 5819 3290 5825 3292
rect 5881 3290 5905 3292
rect 5961 3290 5985 3292
rect 6041 3290 6065 3292
rect 6121 3290 6127 3292
rect 5881 3238 5883 3290
rect 6063 3238 6065 3290
rect 5819 3236 5825 3238
rect 5881 3236 5905 3238
rect 5961 3236 5985 3238
rect 6041 3236 6065 3238
rect 6121 3236 6127 3238
rect 5819 3227 6127 3236
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 6196 2854 6224 3454
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 3194 6316 3334
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6840 2990 6868 3470
rect 6932 3194 6960 3674
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7024 3058 7052 5646
rect 7208 3194 7236 6666
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 5778 7328 6598
rect 8312 6458 8340 6734
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 7965 6012 8273 6021
rect 7965 6010 7971 6012
rect 8027 6010 8051 6012
rect 8107 6010 8131 6012
rect 8187 6010 8211 6012
rect 8267 6010 8273 6012
rect 8027 5958 8029 6010
rect 8209 5958 8211 6010
rect 7965 5956 7971 5958
rect 8027 5956 8051 5958
rect 8107 5956 8131 5958
rect 8187 5956 8211 5958
rect 8267 5956 8273 5958
rect 7965 5947 8273 5956
rect 8404 5914 8432 6854
rect 8772 6798 8800 6870
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8625 6556 8933 6565
rect 8625 6554 8631 6556
rect 8687 6554 8711 6556
rect 8767 6554 8791 6556
rect 8847 6554 8871 6556
rect 8927 6554 8933 6556
rect 8687 6502 8689 6554
rect 8869 6502 8871 6554
rect 8625 6500 8631 6502
rect 8687 6500 8711 6502
rect 8767 6500 8791 6502
rect 8847 6500 8871 6502
rect 8927 6500 8933 6502
rect 8625 6491 8933 6500
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8680 5914 8708 6258
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8312 5370 8340 5578
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 3602 7328 4082
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7300 3126 7328 3334
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6196 2650 6224 2790
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6840 2446 6868 2926
rect 7392 2514 7420 5102
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7576 4146 7604 4490
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3534 7512 3878
rect 7576 3534 7604 3946
rect 7668 3738 7696 4082
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7760 3398 7788 5238
rect 7965 4924 8273 4933
rect 7965 4922 7971 4924
rect 8027 4922 8051 4924
rect 8107 4922 8131 4924
rect 8187 4922 8211 4924
rect 8267 4922 8273 4924
rect 8027 4870 8029 4922
rect 8209 4870 8211 4922
rect 7965 4868 7971 4870
rect 8027 4868 8051 4870
rect 8107 4868 8131 4870
rect 8187 4868 8211 4870
rect 8267 4868 8273 4870
rect 7965 4859 8273 4868
rect 8404 4758 8432 5850
rect 8625 5468 8933 5477
rect 8625 5466 8631 5468
rect 8687 5466 8711 5468
rect 8767 5466 8791 5468
rect 8847 5466 8871 5468
rect 8927 5466 8933 5468
rect 8687 5414 8689 5466
rect 8869 5414 8871 5466
rect 8625 5412 8631 5414
rect 8687 5412 8711 5414
rect 8767 5412 8791 5414
rect 8847 5412 8871 5414
rect 8927 5412 8933 5414
rect 8625 5403 8933 5412
rect 9048 4826 9076 8502
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9140 7546 9168 7754
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9600 7410 9628 10474
rect 9876 10130 9904 10610
rect 10152 10606 10180 11698
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10428 10742 10456 11290
rect 10704 10810 10732 11698
rect 10771 11452 11079 11461
rect 10771 11450 10777 11452
rect 10833 11450 10857 11452
rect 10913 11450 10937 11452
rect 10993 11450 11017 11452
rect 11073 11450 11079 11452
rect 10833 11398 10835 11450
rect 11015 11398 11017 11450
rect 10771 11396 10777 11398
rect 10833 11396 10857 11398
rect 10913 11396 10937 11398
rect 10993 11396 11017 11398
rect 11073 11396 11079 11398
rect 10771 11387 11079 11396
rect 11164 11150 11192 11698
rect 11256 11354 11284 12174
rect 11431 11996 11739 12005
rect 11431 11994 11437 11996
rect 11493 11994 11517 11996
rect 11573 11994 11597 11996
rect 11653 11994 11677 11996
rect 11733 11994 11739 11996
rect 11493 11942 11495 11994
rect 11675 11942 11677 11994
rect 11431 11940 11437 11942
rect 11493 11940 11517 11942
rect 11573 11940 11597 11942
rect 11653 11940 11677 11942
rect 11733 11940 11739 11942
rect 11431 11931 11739 11940
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11348 11286 11376 11630
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10152 10266 10180 10542
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9876 9722 9904 10066
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8498 10180 8910
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10060 7546 10088 8434
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10428 8090 10456 8366
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10520 7886 10548 9114
rect 10704 9110 10732 10746
rect 10796 10674 10824 11086
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10888 10606 10916 11086
rect 10980 10810 11008 11086
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11164 10674 11192 11086
rect 11348 10674 11376 11222
rect 11431 10908 11739 10917
rect 11431 10906 11437 10908
rect 11493 10906 11517 10908
rect 11573 10906 11597 10908
rect 11653 10906 11677 10908
rect 11733 10906 11739 10908
rect 11493 10854 11495 10906
rect 11675 10854 11677 10906
rect 11431 10852 11437 10854
rect 11493 10852 11517 10854
rect 11573 10852 11597 10854
rect 11653 10852 11677 10854
rect 11733 10852 11739 10854
rect 11431 10843 11739 10852
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10771 10364 11079 10373
rect 10771 10362 10777 10364
rect 10833 10362 10857 10364
rect 10913 10362 10937 10364
rect 10993 10362 11017 10364
rect 11073 10362 11079 10364
rect 10833 10310 10835 10362
rect 11015 10310 11017 10362
rect 10771 10308 10777 10310
rect 10833 10308 10857 10310
rect 10913 10308 10937 10310
rect 10993 10308 11017 10310
rect 11073 10308 11079 10310
rect 10771 10299 11079 10308
rect 10771 9276 11079 9285
rect 10771 9274 10777 9276
rect 10833 9274 10857 9276
rect 10913 9274 10937 9276
rect 10993 9274 11017 9276
rect 11073 9274 11079 9276
rect 10833 9222 10835 9274
rect 11015 9222 11017 9274
rect 10771 9220 10777 9222
rect 10833 9220 10857 9222
rect 10913 9220 10937 9222
rect 10993 9220 11017 9222
rect 11073 9220 11079 9222
rect 10771 9211 11079 9220
rect 10692 9104 10744 9110
rect 11164 9058 11192 10610
rect 11348 9450 11376 10610
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11431 9820 11739 9829
rect 11431 9818 11437 9820
rect 11493 9818 11517 9820
rect 11573 9818 11597 9820
rect 11653 9818 11677 9820
rect 11733 9818 11739 9820
rect 11493 9766 11495 9818
rect 11675 9766 11677 9818
rect 11431 9764 11437 9766
rect 11493 9764 11517 9766
rect 11573 9764 11597 9766
rect 11653 9764 11677 9766
rect 11733 9764 11739 9766
rect 11431 9755 11739 9764
rect 11992 9625 12020 9998
rect 11978 9616 12034 9625
rect 11978 9551 12034 9560
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 10692 9046 10744 9052
rect 11072 9030 11192 9058
rect 11072 8566 11100 9030
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11886 8936 11942 8945
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 10771 8188 11079 8197
rect 10771 8186 10777 8188
rect 10833 8186 10857 8188
rect 10913 8186 10937 8188
rect 10993 8186 11017 8188
rect 11073 8186 11079 8188
rect 10833 8134 10835 8186
rect 11015 8134 11017 8186
rect 10771 8132 10777 8134
rect 10833 8132 10857 8134
rect 10913 8132 10937 8134
rect 10993 8132 11017 8134
rect 11073 8132 11079 8134
rect 10771 8123 11079 8132
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 4826 9628 7142
rect 9784 7002 9812 7278
rect 10336 7002 10364 7822
rect 10520 7546 10548 7822
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 9692 6798 9720 6938
rect 10428 6934 10456 7278
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9784 6730 9812 6802
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9968 6662 9996 6870
rect 10520 6798 10548 7346
rect 10704 7290 10732 7346
rect 10612 7262 10732 7290
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10612 6746 10640 7262
rect 10796 7188 10824 7346
rect 10704 7160 10824 7188
rect 10704 7002 10732 7160
rect 10771 7100 11079 7109
rect 10771 7098 10777 7100
rect 10833 7098 10857 7100
rect 10913 7098 10937 7100
rect 10993 7098 11017 7100
rect 11073 7098 11079 7100
rect 10833 7046 10835 7098
rect 11015 7046 11017 7098
rect 10771 7044 10777 7046
rect 10833 7044 10857 7046
rect 10913 7044 10937 7046
rect 10993 7044 11017 7046
rect 11073 7044 11079 7046
rect 10771 7035 11079 7044
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10692 6792 10744 6798
rect 10612 6740 10692 6746
rect 10612 6734 10744 6740
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4146 8340 4422
rect 8404 4282 8432 4694
rect 9048 4622 9076 4762
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 8625 4380 8933 4389
rect 8625 4378 8631 4380
rect 8687 4378 8711 4380
rect 8767 4378 8791 4380
rect 8847 4378 8871 4380
rect 8927 4378 8933 4380
rect 8687 4326 8689 4378
rect 8869 4326 8871 4378
rect 8625 4324 8631 4326
rect 8687 4324 8711 4326
rect 8767 4324 8791 4326
rect 8847 4324 8871 4326
rect 8927 4324 8933 4326
rect 8625 4315 8933 4324
rect 9324 4282 9352 4422
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7852 3534 7880 4014
rect 7965 3836 8273 3845
rect 7965 3834 7971 3836
rect 8027 3834 8051 3836
rect 8107 3834 8131 3836
rect 8187 3834 8211 3836
rect 8267 3834 8273 3836
rect 8027 3782 8029 3834
rect 8209 3782 8211 3834
rect 7965 3780 7971 3782
rect 8027 3780 8051 3782
rect 8107 3780 8131 3782
rect 8187 3780 8211 3782
rect 8267 3780 8273 3782
rect 7965 3771 8273 3780
rect 8956 3738 8984 4082
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7852 2774 7880 3470
rect 7944 3194 7972 3674
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8036 3126 8064 3334
rect 8625 3292 8933 3301
rect 8625 3290 8631 3292
rect 8687 3290 8711 3292
rect 8767 3290 8791 3292
rect 8847 3290 8871 3292
rect 8927 3290 8933 3292
rect 8687 3238 8689 3290
rect 8869 3238 8871 3290
rect 8625 3236 8631 3238
rect 8687 3236 8711 3238
rect 8767 3236 8791 3238
rect 8847 3236 8871 3238
rect 8927 3236 8933 3238
rect 8625 3227 8933 3236
rect 9048 3194 9076 4150
rect 9692 3738 9720 4422
rect 9968 4146 9996 6598
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5846 10088 6258
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10060 4622 10088 5782
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10152 4554 10180 6734
rect 10612 6718 10732 6734
rect 10704 6458 10732 6718
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10888 6322 10916 6870
rect 11164 6662 11192 8910
rect 11886 8871 11942 8880
rect 11431 8732 11739 8741
rect 11431 8730 11437 8732
rect 11493 8730 11517 8732
rect 11573 8730 11597 8732
rect 11653 8730 11677 8732
rect 11733 8730 11739 8732
rect 11493 8678 11495 8730
rect 11675 8678 11677 8730
rect 11431 8676 11437 8678
rect 11493 8676 11517 8678
rect 11573 8676 11597 8678
rect 11653 8676 11677 8678
rect 11733 8676 11739 8678
rect 11431 8667 11739 8676
rect 11900 8634 11928 8871
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11431 7644 11739 7653
rect 11431 7642 11437 7644
rect 11493 7642 11517 7644
rect 11573 7642 11597 7644
rect 11653 7642 11677 7644
rect 11733 7642 11739 7644
rect 11493 7590 11495 7642
rect 11675 7590 11677 7642
rect 11431 7588 11437 7590
rect 11493 7588 11517 7590
rect 11573 7588 11597 7590
rect 11653 7588 11677 7590
rect 11733 7588 11739 7590
rect 11431 7579 11739 7588
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6458 11192 6598
rect 11256 6458 11284 6666
rect 11431 6556 11739 6565
rect 11431 6554 11437 6556
rect 11493 6554 11517 6556
rect 11573 6554 11597 6556
rect 11653 6554 11677 6556
rect 11733 6554 11739 6556
rect 11493 6502 11495 6554
rect 11675 6502 11677 6554
rect 11431 6500 11437 6502
rect 11493 6500 11517 6502
rect 11573 6500 11597 6502
rect 11653 6500 11677 6502
rect 11733 6500 11739 6502
rect 11431 6491 11739 6500
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 10704 5914 10732 6258
rect 10771 6012 11079 6021
rect 10771 6010 10777 6012
rect 10833 6010 10857 6012
rect 10913 6010 10937 6012
rect 10993 6010 11017 6012
rect 11073 6010 11079 6012
rect 10833 5958 10835 6010
rect 11015 5958 11017 6010
rect 10771 5956 10777 5958
rect 10833 5956 10857 5958
rect 10913 5956 10937 5958
rect 10993 5956 11017 5958
rect 11073 5956 11079 5958
rect 10771 5947 11079 5956
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 11348 5846 11376 6258
rect 11886 6216 11942 6225
rect 11886 6151 11888 6160
rect 11940 6151 11942 6160
rect 11888 6122 11940 6128
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 10520 5166 10548 5646
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9416 3194 9444 3470
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9692 3126 9720 3674
rect 9784 3670 9812 4082
rect 9968 4010 9996 4082
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 10152 3738 10180 4490
rect 10244 4214 10272 4626
rect 10520 4622 10548 5102
rect 10704 5030 10732 5646
rect 11992 5545 12020 5646
rect 11978 5536 12034 5545
rect 11431 5468 11739 5477
rect 11978 5471 12034 5480
rect 11431 5466 11437 5468
rect 11493 5466 11517 5468
rect 11573 5466 11597 5468
rect 11653 5466 11677 5468
rect 11733 5466 11739 5468
rect 11493 5414 11495 5466
rect 11675 5414 11677 5466
rect 11431 5412 11437 5414
rect 11493 5412 11517 5414
rect 11573 5412 11597 5414
rect 11653 5412 11677 5414
rect 11733 5412 11739 5414
rect 11431 5403 11739 5412
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4758 10732 4966
rect 10771 4924 11079 4933
rect 10771 4922 10777 4924
rect 10833 4922 10857 4924
rect 10913 4922 10937 4924
rect 10993 4922 11017 4924
rect 11073 4922 11079 4924
rect 10833 4870 10835 4922
rect 11015 4870 11017 4922
rect 10771 4868 10777 4870
rect 10833 4868 10857 4870
rect 10913 4868 10937 4870
rect 10993 4868 11017 4870
rect 11073 4868 11079 4870
rect 10771 4859 11079 4868
rect 11992 4865 12020 5170
rect 11978 4856 12034 4865
rect 11978 4791 12034 4800
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10704 4622 10732 4694
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 11256 4146 11284 4490
rect 11431 4380 11739 4389
rect 11431 4378 11437 4380
rect 11493 4378 11517 4380
rect 11573 4378 11597 4380
rect 11653 4378 11677 4380
rect 11733 4378 11739 4380
rect 11493 4326 11495 4378
rect 11675 4326 11677 4378
rect 11431 4324 11437 4326
rect 11493 4324 11517 4326
rect 11573 4324 11597 4326
rect 11653 4324 11677 4326
rect 11733 4324 11739 4326
rect 11431 4315 11739 4324
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 10244 3534 10272 3946
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9692 2854 9720 3062
rect 9784 3058 9812 3470
rect 10428 3058 10456 4014
rect 10612 3942 10640 4082
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 10612 3670 10640 3878
rect 10771 3836 11079 3845
rect 10771 3834 10777 3836
rect 10833 3834 10857 3836
rect 10913 3834 10937 3836
rect 10993 3834 11017 3836
rect 11073 3834 11079 3836
rect 10833 3782 10835 3834
rect 11015 3782 11017 3834
rect 10771 3780 10777 3782
rect 10833 3780 10857 3782
rect 10913 3780 10937 3782
rect 10993 3780 11017 3782
rect 11073 3780 11079 3782
rect 10771 3771 11079 3780
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10612 2990 10640 3606
rect 11624 3534 11652 3878
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11886 3496 11942 3505
rect 11886 3431 11888 3440
rect 11940 3431 11942 3440
rect 11888 3402 11940 3408
rect 11431 3292 11739 3301
rect 11431 3290 11437 3292
rect 11493 3290 11517 3292
rect 11573 3290 11597 3292
rect 11653 3290 11677 3292
rect 11733 3290 11739 3292
rect 11493 3238 11495 3290
rect 11675 3238 11677 3290
rect 11431 3236 11437 3238
rect 11493 3236 11517 3238
rect 11573 3236 11597 3238
rect 11653 3236 11677 3238
rect 11733 3236 11739 3238
rect 11431 3227 11739 3236
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 7668 2746 7880 2774
rect 7965 2748 8273 2757
rect 7965 2746 7971 2748
rect 8027 2746 8051 2748
rect 8107 2746 8131 2748
rect 8187 2746 8211 2748
rect 8267 2746 8273 2748
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7668 2446 7696 2746
rect 8027 2694 8029 2746
rect 8209 2694 8211 2746
rect 7965 2692 7971 2694
rect 8027 2692 8051 2694
rect 8107 2692 8131 2694
rect 8187 2692 8211 2694
rect 8267 2692 8273 2694
rect 7965 2683 8273 2692
rect 10771 2748 11079 2757
rect 10771 2746 10777 2748
rect 10833 2746 10857 2748
rect 10913 2746 10937 2748
rect 10993 2746 11017 2748
rect 11073 2746 11079 2748
rect 10833 2694 10835 2746
rect 11015 2694 11017 2746
rect 10771 2692 10777 2694
rect 10833 2692 10857 2694
rect 10913 2692 10937 2694
rect 10993 2692 11017 2694
rect 11073 2692 11079 2694
rect 10771 2683 11079 2692
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 3013 2204 3321 2213
rect 3013 2202 3019 2204
rect 3075 2202 3099 2204
rect 3155 2202 3179 2204
rect 3235 2202 3259 2204
rect 3315 2202 3321 2204
rect 3075 2150 3077 2202
rect 3257 2150 3259 2202
rect 3013 2148 3019 2150
rect 3075 2148 3099 2150
rect 3155 2148 3179 2150
rect 3235 2148 3259 2150
rect 3315 2148 3321 2150
rect 3013 2139 3321 2148
rect 5736 1306 5764 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 5819 2204 6127 2213
rect 5819 2202 5825 2204
rect 5881 2202 5905 2204
rect 5961 2202 5985 2204
rect 6041 2202 6065 2204
rect 6121 2202 6127 2204
rect 5881 2150 5883 2202
rect 6063 2150 6065 2202
rect 5819 2148 5825 2150
rect 5881 2148 5905 2150
rect 5961 2148 5985 2150
rect 6041 2148 6065 2150
rect 6121 2148 6127 2150
rect 5819 2139 6127 2148
rect 5736 1278 5856 1306
rect 5828 800 5856 1278
rect 6472 800 6500 2246
rect 7116 800 7144 2246
rect 7760 800 7788 2246
rect 8625 2204 8933 2213
rect 8625 2202 8631 2204
rect 8687 2202 8711 2204
rect 8767 2202 8791 2204
rect 8847 2202 8871 2204
rect 8927 2202 8933 2204
rect 8687 2150 8689 2202
rect 8869 2150 8871 2202
rect 8625 2148 8631 2150
rect 8687 2148 8711 2150
rect 8767 2148 8791 2150
rect 8847 2148 8871 2150
rect 8927 2148 8933 2150
rect 8625 2139 8933 2148
rect 11431 2204 11739 2213
rect 11431 2202 11437 2204
rect 11493 2202 11517 2204
rect 11573 2202 11597 2204
rect 11653 2202 11677 2204
rect 11733 2202 11739 2204
rect 11493 2150 11495 2202
rect 11675 2150 11677 2202
rect 11431 2148 11437 2150
rect 11493 2148 11517 2150
rect 11573 2148 11597 2150
rect 11653 2148 11677 2150
rect 11733 2148 11739 2150
rect 11431 2139 11739 2148
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
<< via2 >>
rect 3019 13082 3075 13084
rect 3099 13082 3155 13084
rect 3179 13082 3235 13084
rect 3259 13082 3315 13084
rect 3019 13030 3065 13082
rect 3065 13030 3075 13082
rect 3099 13030 3129 13082
rect 3129 13030 3141 13082
rect 3141 13030 3155 13082
rect 3179 13030 3193 13082
rect 3193 13030 3205 13082
rect 3205 13030 3235 13082
rect 3259 13030 3269 13082
rect 3269 13030 3315 13082
rect 3019 13028 3075 13030
rect 3099 13028 3155 13030
rect 3179 13028 3235 13030
rect 3259 13028 3315 13030
rect 5825 13082 5881 13084
rect 5905 13082 5961 13084
rect 5985 13082 6041 13084
rect 6065 13082 6121 13084
rect 5825 13030 5871 13082
rect 5871 13030 5881 13082
rect 5905 13030 5935 13082
rect 5935 13030 5947 13082
rect 5947 13030 5961 13082
rect 5985 13030 5999 13082
rect 5999 13030 6011 13082
rect 6011 13030 6041 13082
rect 6065 13030 6075 13082
rect 6075 13030 6121 13082
rect 5825 13028 5881 13030
rect 5905 13028 5961 13030
rect 5985 13028 6041 13030
rect 6065 13028 6121 13030
rect 8631 13082 8687 13084
rect 8711 13082 8767 13084
rect 8791 13082 8847 13084
rect 8871 13082 8927 13084
rect 8631 13030 8677 13082
rect 8677 13030 8687 13082
rect 8711 13030 8741 13082
rect 8741 13030 8753 13082
rect 8753 13030 8767 13082
rect 8791 13030 8805 13082
rect 8805 13030 8817 13082
rect 8817 13030 8847 13082
rect 8871 13030 8881 13082
rect 8881 13030 8927 13082
rect 8631 13028 8687 13030
rect 8711 13028 8767 13030
rect 8791 13028 8847 13030
rect 8871 13028 8927 13030
rect 11437 13082 11493 13084
rect 11517 13082 11573 13084
rect 11597 13082 11653 13084
rect 11677 13082 11733 13084
rect 11437 13030 11483 13082
rect 11483 13030 11493 13082
rect 11517 13030 11547 13082
rect 11547 13030 11559 13082
rect 11559 13030 11573 13082
rect 11597 13030 11611 13082
rect 11611 13030 11623 13082
rect 11623 13030 11653 13082
rect 11677 13030 11687 13082
rect 11687 13030 11733 13082
rect 11437 13028 11493 13030
rect 11517 13028 11573 13030
rect 11597 13028 11653 13030
rect 11677 13028 11733 13030
rect 2359 12538 2415 12540
rect 2439 12538 2495 12540
rect 2519 12538 2575 12540
rect 2599 12538 2655 12540
rect 2359 12486 2405 12538
rect 2405 12486 2415 12538
rect 2439 12486 2469 12538
rect 2469 12486 2481 12538
rect 2481 12486 2495 12538
rect 2519 12486 2533 12538
rect 2533 12486 2545 12538
rect 2545 12486 2575 12538
rect 2599 12486 2609 12538
rect 2609 12486 2655 12538
rect 2359 12484 2415 12486
rect 2439 12484 2495 12486
rect 2519 12484 2575 12486
rect 2599 12484 2655 12486
rect 5165 12538 5221 12540
rect 5245 12538 5301 12540
rect 5325 12538 5381 12540
rect 5405 12538 5461 12540
rect 5165 12486 5211 12538
rect 5211 12486 5221 12538
rect 5245 12486 5275 12538
rect 5275 12486 5287 12538
rect 5287 12486 5301 12538
rect 5325 12486 5339 12538
rect 5339 12486 5351 12538
rect 5351 12486 5381 12538
rect 5405 12486 5415 12538
rect 5415 12486 5461 12538
rect 5165 12484 5221 12486
rect 5245 12484 5301 12486
rect 5325 12484 5381 12486
rect 5405 12484 5461 12486
rect 3019 11994 3075 11996
rect 3099 11994 3155 11996
rect 3179 11994 3235 11996
rect 3259 11994 3315 11996
rect 3019 11942 3065 11994
rect 3065 11942 3075 11994
rect 3099 11942 3129 11994
rect 3129 11942 3141 11994
rect 3141 11942 3155 11994
rect 3179 11942 3193 11994
rect 3193 11942 3205 11994
rect 3205 11942 3235 11994
rect 3259 11942 3269 11994
rect 3269 11942 3315 11994
rect 3019 11940 3075 11942
rect 3099 11940 3155 11942
rect 3179 11940 3235 11942
rect 3259 11940 3315 11942
rect 2359 11450 2415 11452
rect 2439 11450 2495 11452
rect 2519 11450 2575 11452
rect 2599 11450 2655 11452
rect 2359 11398 2405 11450
rect 2405 11398 2415 11450
rect 2439 11398 2469 11450
rect 2469 11398 2481 11450
rect 2481 11398 2495 11450
rect 2519 11398 2533 11450
rect 2533 11398 2545 11450
rect 2545 11398 2575 11450
rect 2599 11398 2609 11450
rect 2609 11398 2655 11450
rect 2359 11396 2415 11398
rect 2439 11396 2495 11398
rect 2519 11396 2575 11398
rect 2599 11396 2655 11398
rect 1398 10920 1454 10976
rect 1306 10260 1362 10296
rect 1306 10240 1308 10260
rect 1308 10240 1360 10260
rect 1360 10240 1362 10260
rect 2359 10362 2415 10364
rect 2439 10362 2495 10364
rect 2519 10362 2575 10364
rect 2599 10362 2655 10364
rect 2359 10310 2405 10362
rect 2405 10310 2415 10362
rect 2439 10310 2469 10362
rect 2469 10310 2481 10362
rect 2481 10310 2495 10362
rect 2519 10310 2533 10362
rect 2533 10310 2545 10362
rect 2545 10310 2575 10362
rect 2599 10310 2609 10362
rect 2609 10310 2655 10362
rect 2359 10308 2415 10310
rect 2439 10308 2495 10310
rect 2519 10308 2575 10310
rect 2599 10308 2655 10310
rect 5825 11994 5881 11996
rect 5905 11994 5961 11996
rect 5985 11994 6041 11996
rect 6065 11994 6121 11996
rect 5825 11942 5871 11994
rect 5871 11942 5881 11994
rect 5905 11942 5935 11994
rect 5935 11942 5947 11994
rect 5947 11942 5961 11994
rect 5985 11942 5999 11994
rect 5999 11942 6011 11994
rect 6011 11942 6041 11994
rect 6065 11942 6075 11994
rect 6075 11942 6121 11994
rect 5825 11940 5881 11942
rect 5905 11940 5961 11942
rect 5985 11940 6041 11942
rect 6065 11940 6121 11942
rect 5165 11450 5221 11452
rect 5245 11450 5301 11452
rect 5325 11450 5381 11452
rect 5405 11450 5461 11452
rect 5165 11398 5211 11450
rect 5211 11398 5221 11450
rect 5245 11398 5275 11450
rect 5275 11398 5287 11450
rect 5287 11398 5301 11450
rect 5325 11398 5339 11450
rect 5339 11398 5351 11450
rect 5351 11398 5381 11450
rect 5405 11398 5415 11450
rect 5415 11398 5461 11450
rect 5165 11396 5221 11398
rect 5245 11396 5301 11398
rect 5325 11396 5381 11398
rect 5405 11396 5461 11398
rect 3019 10906 3075 10908
rect 3099 10906 3155 10908
rect 3179 10906 3235 10908
rect 3259 10906 3315 10908
rect 3019 10854 3065 10906
rect 3065 10854 3075 10906
rect 3099 10854 3129 10906
rect 3129 10854 3141 10906
rect 3141 10854 3155 10906
rect 3179 10854 3193 10906
rect 3193 10854 3205 10906
rect 3205 10854 3235 10906
rect 3259 10854 3269 10906
rect 3269 10854 3315 10906
rect 3019 10852 3075 10854
rect 3099 10852 3155 10854
rect 3179 10852 3235 10854
rect 3259 10852 3315 10854
rect 3019 9818 3075 9820
rect 3099 9818 3155 9820
rect 3179 9818 3235 9820
rect 3259 9818 3315 9820
rect 3019 9766 3065 9818
rect 3065 9766 3075 9818
rect 3099 9766 3129 9818
rect 3129 9766 3141 9818
rect 3141 9766 3155 9818
rect 3179 9766 3193 9818
rect 3193 9766 3205 9818
rect 3205 9766 3235 9818
rect 3259 9766 3269 9818
rect 3269 9766 3315 9818
rect 3019 9764 3075 9766
rect 3099 9764 3155 9766
rect 3179 9764 3235 9766
rect 3259 9764 3315 9766
rect 2359 9274 2415 9276
rect 2439 9274 2495 9276
rect 2519 9274 2575 9276
rect 2599 9274 2655 9276
rect 2359 9222 2405 9274
rect 2405 9222 2415 9274
rect 2439 9222 2469 9274
rect 2469 9222 2481 9274
rect 2481 9222 2495 9274
rect 2519 9222 2533 9274
rect 2533 9222 2545 9274
rect 2545 9222 2575 9274
rect 2599 9222 2609 9274
rect 2609 9222 2655 9274
rect 2359 9220 2415 9222
rect 2439 9220 2495 9222
rect 2519 9220 2575 9222
rect 2599 9220 2655 9222
rect 5165 10362 5221 10364
rect 5245 10362 5301 10364
rect 5325 10362 5381 10364
rect 5405 10362 5461 10364
rect 5165 10310 5211 10362
rect 5211 10310 5221 10362
rect 5245 10310 5275 10362
rect 5275 10310 5287 10362
rect 5287 10310 5301 10362
rect 5325 10310 5339 10362
rect 5339 10310 5351 10362
rect 5351 10310 5381 10362
rect 5405 10310 5415 10362
rect 5415 10310 5461 10362
rect 5165 10308 5221 10310
rect 5245 10308 5301 10310
rect 5325 10308 5381 10310
rect 5405 10308 5461 10310
rect 3019 8730 3075 8732
rect 3099 8730 3155 8732
rect 3179 8730 3235 8732
rect 3259 8730 3315 8732
rect 3019 8678 3065 8730
rect 3065 8678 3075 8730
rect 3099 8678 3129 8730
rect 3129 8678 3141 8730
rect 3141 8678 3155 8730
rect 3179 8678 3193 8730
rect 3193 8678 3205 8730
rect 3205 8678 3235 8730
rect 3259 8678 3269 8730
rect 3269 8678 3315 8730
rect 3019 8676 3075 8678
rect 3099 8676 3155 8678
rect 3179 8676 3235 8678
rect 3259 8676 3315 8678
rect 1306 8200 1362 8256
rect 2359 8186 2415 8188
rect 2439 8186 2495 8188
rect 2519 8186 2575 8188
rect 2599 8186 2655 8188
rect 2359 8134 2405 8186
rect 2405 8134 2415 8186
rect 2439 8134 2469 8186
rect 2469 8134 2481 8186
rect 2481 8134 2495 8186
rect 2519 8134 2533 8186
rect 2533 8134 2545 8186
rect 2545 8134 2575 8186
rect 2599 8134 2609 8186
rect 2609 8134 2655 8186
rect 2359 8132 2415 8134
rect 2439 8132 2495 8134
rect 2519 8132 2575 8134
rect 2599 8132 2655 8134
rect 2359 7098 2415 7100
rect 2439 7098 2495 7100
rect 2519 7098 2575 7100
rect 2599 7098 2655 7100
rect 2359 7046 2405 7098
rect 2405 7046 2415 7098
rect 2439 7046 2469 7098
rect 2469 7046 2481 7098
rect 2481 7046 2495 7098
rect 2519 7046 2533 7098
rect 2533 7046 2545 7098
rect 2545 7046 2575 7098
rect 2599 7046 2609 7098
rect 2609 7046 2655 7098
rect 2359 7044 2415 7046
rect 2439 7044 2495 7046
rect 2519 7044 2575 7046
rect 2599 7044 2655 7046
rect 2359 6010 2415 6012
rect 2439 6010 2495 6012
rect 2519 6010 2575 6012
rect 2599 6010 2655 6012
rect 2359 5958 2405 6010
rect 2405 5958 2415 6010
rect 2439 5958 2469 6010
rect 2469 5958 2481 6010
rect 2481 5958 2495 6010
rect 2519 5958 2533 6010
rect 2533 5958 2545 6010
rect 2545 5958 2575 6010
rect 2599 5958 2609 6010
rect 2609 5958 2655 6010
rect 2359 5956 2415 5958
rect 2439 5956 2495 5958
rect 2519 5956 2575 5958
rect 2599 5956 2655 5958
rect 2359 4922 2415 4924
rect 2439 4922 2495 4924
rect 2519 4922 2575 4924
rect 2599 4922 2655 4924
rect 2359 4870 2405 4922
rect 2405 4870 2415 4922
rect 2439 4870 2469 4922
rect 2469 4870 2481 4922
rect 2481 4870 2495 4922
rect 2519 4870 2533 4922
rect 2533 4870 2545 4922
rect 2545 4870 2575 4922
rect 2599 4870 2609 4922
rect 2609 4870 2655 4922
rect 2359 4868 2415 4870
rect 2439 4868 2495 4870
rect 2519 4868 2575 4870
rect 2599 4868 2655 4870
rect 3019 7642 3075 7644
rect 3099 7642 3155 7644
rect 3179 7642 3235 7644
rect 3259 7642 3315 7644
rect 3019 7590 3065 7642
rect 3065 7590 3075 7642
rect 3099 7590 3129 7642
rect 3129 7590 3141 7642
rect 3141 7590 3155 7642
rect 3179 7590 3193 7642
rect 3193 7590 3205 7642
rect 3205 7590 3235 7642
rect 3259 7590 3269 7642
rect 3269 7590 3315 7642
rect 3019 7588 3075 7590
rect 3099 7588 3155 7590
rect 3179 7588 3235 7590
rect 3259 7588 3315 7590
rect 3019 6554 3075 6556
rect 3099 6554 3155 6556
rect 3179 6554 3235 6556
rect 3259 6554 3315 6556
rect 3019 6502 3065 6554
rect 3065 6502 3075 6554
rect 3099 6502 3129 6554
rect 3129 6502 3141 6554
rect 3141 6502 3155 6554
rect 3179 6502 3193 6554
rect 3193 6502 3205 6554
rect 3205 6502 3235 6554
rect 3259 6502 3269 6554
rect 3269 6502 3315 6554
rect 3019 6500 3075 6502
rect 3099 6500 3155 6502
rect 3179 6500 3235 6502
rect 3259 6500 3315 6502
rect 3019 5466 3075 5468
rect 3099 5466 3155 5468
rect 3179 5466 3235 5468
rect 3259 5466 3315 5468
rect 3019 5414 3065 5466
rect 3065 5414 3075 5466
rect 3099 5414 3129 5466
rect 3129 5414 3141 5466
rect 3141 5414 3155 5466
rect 3179 5414 3193 5466
rect 3193 5414 3205 5466
rect 3205 5414 3235 5466
rect 3259 5414 3269 5466
rect 3269 5414 3315 5466
rect 3019 5412 3075 5414
rect 3099 5412 3155 5414
rect 3179 5412 3235 5414
rect 3259 5412 3315 5414
rect 4250 8200 4306 8256
rect 5165 9274 5221 9276
rect 5245 9274 5301 9276
rect 5325 9274 5381 9276
rect 5405 9274 5461 9276
rect 5165 9222 5211 9274
rect 5211 9222 5221 9274
rect 5245 9222 5275 9274
rect 5275 9222 5287 9274
rect 5287 9222 5301 9274
rect 5325 9222 5339 9274
rect 5339 9222 5351 9274
rect 5351 9222 5381 9274
rect 5405 9222 5415 9274
rect 5415 9222 5461 9274
rect 5165 9220 5221 9222
rect 5245 9220 5301 9222
rect 5325 9220 5381 9222
rect 5405 9220 5461 9222
rect 5825 10906 5881 10908
rect 5905 10906 5961 10908
rect 5985 10906 6041 10908
rect 6065 10906 6121 10908
rect 5825 10854 5871 10906
rect 5871 10854 5881 10906
rect 5905 10854 5935 10906
rect 5935 10854 5947 10906
rect 5947 10854 5961 10906
rect 5985 10854 5999 10906
rect 5999 10854 6011 10906
rect 6011 10854 6041 10906
rect 6065 10854 6075 10906
rect 6075 10854 6121 10906
rect 5825 10852 5881 10854
rect 5905 10852 5961 10854
rect 5985 10852 6041 10854
rect 6065 10852 6121 10854
rect 5825 9818 5881 9820
rect 5905 9818 5961 9820
rect 5985 9818 6041 9820
rect 6065 9818 6121 9820
rect 5825 9766 5871 9818
rect 5871 9766 5881 9818
rect 5905 9766 5935 9818
rect 5935 9766 5947 9818
rect 5947 9766 5961 9818
rect 5985 9766 5999 9818
rect 5999 9766 6011 9818
rect 6011 9766 6041 9818
rect 6065 9766 6075 9818
rect 6075 9766 6121 9818
rect 5825 9764 5881 9766
rect 5905 9764 5961 9766
rect 5985 9764 6041 9766
rect 6065 9764 6121 9766
rect 5825 8730 5881 8732
rect 5905 8730 5961 8732
rect 5985 8730 6041 8732
rect 6065 8730 6121 8732
rect 5825 8678 5871 8730
rect 5871 8678 5881 8730
rect 5905 8678 5935 8730
rect 5935 8678 5947 8730
rect 5947 8678 5961 8730
rect 5985 8678 5999 8730
rect 5999 8678 6011 8730
rect 6011 8678 6041 8730
rect 6065 8678 6075 8730
rect 6075 8678 6121 8730
rect 5825 8676 5881 8678
rect 5905 8676 5961 8678
rect 5985 8676 6041 8678
rect 6065 8676 6121 8678
rect 5165 8186 5221 8188
rect 5245 8186 5301 8188
rect 5325 8186 5381 8188
rect 5405 8186 5461 8188
rect 5165 8134 5211 8186
rect 5211 8134 5221 8186
rect 5245 8134 5275 8186
rect 5275 8134 5287 8186
rect 5287 8134 5301 8186
rect 5325 8134 5339 8186
rect 5339 8134 5351 8186
rect 5351 8134 5381 8186
rect 5405 8134 5415 8186
rect 5415 8134 5461 8186
rect 5165 8132 5221 8134
rect 5245 8132 5301 8134
rect 5325 8132 5381 8134
rect 5405 8132 5461 8134
rect 7971 12538 8027 12540
rect 8051 12538 8107 12540
rect 8131 12538 8187 12540
rect 8211 12538 8267 12540
rect 7971 12486 8017 12538
rect 8017 12486 8027 12538
rect 8051 12486 8081 12538
rect 8081 12486 8093 12538
rect 8093 12486 8107 12538
rect 8131 12486 8145 12538
rect 8145 12486 8157 12538
rect 8157 12486 8187 12538
rect 8211 12486 8221 12538
rect 8221 12486 8267 12538
rect 7971 12484 8027 12486
rect 8051 12484 8107 12486
rect 8131 12484 8187 12486
rect 8211 12484 8267 12486
rect 7971 11450 8027 11452
rect 8051 11450 8107 11452
rect 8131 11450 8187 11452
rect 8211 11450 8267 11452
rect 7971 11398 8017 11450
rect 8017 11398 8027 11450
rect 8051 11398 8081 11450
rect 8081 11398 8093 11450
rect 8093 11398 8107 11450
rect 8131 11398 8145 11450
rect 8145 11398 8157 11450
rect 8157 11398 8187 11450
rect 8211 11398 8221 11450
rect 8221 11398 8267 11450
rect 7971 11396 8027 11398
rect 8051 11396 8107 11398
rect 8131 11396 8187 11398
rect 8211 11396 8267 11398
rect 7971 10362 8027 10364
rect 8051 10362 8107 10364
rect 8131 10362 8187 10364
rect 8211 10362 8267 10364
rect 7971 10310 8017 10362
rect 8017 10310 8027 10362
rect 8051 10310 8081 10362
rect 8081 10310 8093 10362
rect 8093 10310 8107 10362
rect 8131 10310 8145 10362
rect 8145 10310 8157 10362
rect 8157 10310 8187 10362
rect 8211 10310 8221 10362
rect 8221 10310 8267 10362
rect 7971 10308 8027 10310
rect 8051 10308 8107 10310
rect 8131 10308 8187 10310
rect 8211 10308 8267 10310
rect 7971 9274 8027 9276
rect 8051 9274 8107 9276
rect 8131 9274 8187 9276
rect 8211 9274 8267 9276
rect 7971 9222 8017 9274
rect 8017 9222 8027 9274
rect 8051 9222 8081 9274
rect 8081 9222 8093 9274
rect 8093 9222 8107 9274
rect 8131 9222 8145 9274
rect 8145 9222 8157 9274
rect 8157 9222 8187 9274
rect 8211 9222 8221 9274
rect 8221 9222 8267 9274
rect 7971 9220 8027 9222
rect 8051 9220 8107 9222
rect 8131 9220 8187 9222
rect 8211 9220 8267 9222
rect 5825 7642 5881 7644
rect 5905 7642 5961 7644
rect 5985 7642 6041 7644
rect 6065 7642 6121 7644
rect 5825 7590 5871 7642
rect 5871 7590 5881 7642
rect 5905 7590 5935 7642
rect 5935 7590 5947 7642
rect 5947 7590 5961 7642
rect 5985 7590 5999 7642
rect 5999 7590 6011 7642
rect 6011 7590 6041 7642
rect 6065 7590 6075 7642
rect 6075 7590 6121 7642
rect 5825 7588 5881 7590
rect 5905 7588 5961 7590
rect 5985 7588 6041 7590
rect 6065 7588 6121 7590
rect 5165 7098 5221 7100
rect 5245 7098 5301 7100
rect 5325 7098 5381 7100
rect 5405 7098 5461 7100
rect 5165 7046 5211 7098
rect 5211 7046 5221 7098
rect 5245 7046 5275 7098
rect 5275 7046 5287 7098
rect 5287 7046 5301 7098
rect 5325 7046 5339 7098
rect 5339 7046 5351 7098
rect 5351 7046 5381 7098
rect 5405 7046 5415 7098
rect 5415 7046 5461 7098
rect 5165 7044 5221 7046
rect 5245 7044 5301 7046
rect 5325 7044 5381 7046
rect 5405 7044 5461 7046
rect 3019 4378 3075 4380
rect 3099 4378 3155 4380
rect 3179 4378 3235 4380
rect 3259 4378 3315 4380
rect 3019 4326 3065 4378
rect 3065 4326 3075 4378
rect 3099 4326 3129 4378
rect 3129 4326 3141 4378
rect 3141 4326 3155 4378
rect 3179 4326 3193 4378
rect 3193 4326 3205 4378
rect 3205 4326 3235 4378
rect 3259 4326 3269 4378
rect 3269 4326 3315 4378
rect 3019 4324 3075 4326
rect 3099 4324 3155 4326
rect 3179 4324 3235 4326
rect 3259 4324 3315 4326
rect 2359 3834 2415 3836
rect 2439 3834 2495 3836
rect 2519 3834 2575 3836
rect 2599 3834 2655 3836
rect 2359 3782 2405 3834
rect 2405 3782 2415 3834
rect 2439 3782 2469 3834
rect 2469 3782 2481 3834
rect 2481 3782 2495 3834
rect 2519 3782 2533 3834
rect 2533 3782 2545 3834
rect 2545 3782 2575 3834
rect 2599 3782 2609 3834
rect 2609 3782 2655 3834
rect 2359 3780 2415 3782
rect 2439 3780 2495 3782
rect 2519 3780 2575 3782
rect 2599 3780 2655 3782
rect 3019 3290 3075 3292
rect 3099 3290 3155 3292
rect 3179 3290 3235 3292
rect 3259 3290 3315 3292
rect 3019 3238 3065 3290
rect 3065 3238 3075 3290
rect 3099 3238 3129 3290
rect 3129 3238 3141 3290
rect 3141 3238 3155 3290
rect 3179 3238 3193 3290
rect 3193 3238 3205 3290
rect 3205 3238 3235 3290
rect 3259 3238 3269 3290
rect 3269 3238 3315 3290
rect 3019 3236 3075 3238
rect 3099 3236 3155 3238
rect 3179 3236 3235 3238
rect 3259 3236 3315 3238
rect 5165 6010 5221 6012
rect 5245 6010 5301 6012
rect 5325 6010 5381 6012
rect 5405 6010 5461 6012
rect 5165 5958 5211 6010
rect 5211 5958 5221 6010
rect 5245 5958 5275 6010
rect 5275 5958 5287 6010
rect 5287 5958 5301 6010
rect 5325 5958 5339 6010
rect 5339 5958 5351 6010
rect 5351 5958 5381 6010
rect 5405 5958 5415 6010
rect 5415 5958 5461 6010
rect 5165 5956 5221 5958
rect 5245 5956 5301 5958
rect 5325 5956 5381 5958
rect 5405 5956 5461 5958
rect 5825 6554 5881 6556
rect 5905 6554 5961 6556
rect 5985 6554 6041 6556
rect 6065 6554 6121 6556
rect 5825 6502 5871 6554
rect 5871 6502 5881 6554
rect 5905 6502 5935 6554
rect 5935 6502 5947 6554
rect 5947 6502 5961 6554
rect 5985 6502 5999 6554
rect 5999 6502 6011 6554
rect 6011 6502 6041 6554
rect 6065 6502 6075 6554
rect 6075 6502 6121 6554
rect 5825 6500 5881 6502
rect 5905 6500 5961 6502
rect 5985 6500 6041 6502
rect 6065 6500 6121 6502
rect 5165 4922 5221 4924
rect 5245 4922 5301 4924
rect 5325 4922 5381 4924
rect 5405 4922 5461 4924
rect 5165 4870 5211 4922
rect 5211 4870 5221 4922
rect 5245 4870 5275 4922
rect 5275 4870 5287 4922
rect 5287 4870 5301 4922
rect 5325 4870 5339 4922
rect 5339 4870 5351 4922
rect 5351 4870 5381 4922
rect 5405 4870 5415 4922
rect 5415 4870 5461 4922
rect 5165 4868 5221 4870
rect 5245 4868 5301 4870
rect 5325 4868 5381 4870
rect 5405 4868 5461 4870
rect 5825 5466 5881 5468
rect 5905 5466 5961 5468
rect 5985 5466 6041 5468
rect 6065 5466 6121 5468
rect 5825 5414 5871 5466
rect 5871 5414 5881 5466
rect 5905 5414 5935 5466
rect 5935 5414 5947 5466
rect 5947 5414 5961 5466
rect 5985 5414 5999 5466
rect 5999 5414 6011 5466
rect 6011 5414 6041 5466
rect 6065 5414 6075 5466
rect 6075 5414 6121 5466
rect 5825 5412 5881 5414
rect 5905 5412 5961 5414
rect 5985 5412 6041 5414
rect 6065 5412 6121 5414
rect 5165 3834 5221 3836
rect 5245 3834 5301 3836
rect 5325 3834 5381 3836
rect 5405 3834 5461 3836
rect 5165 3782 5211 3834
rect 5211 3782 5221 3834
rect 5245 3782 5275 3834
rect 5275 3782 5287 3834
rect 5287 3782 5301 3834
rect 5325 3782 5339 3834
rect 5339 3782 5351 3834
rect 5351 3782 5381 3834
rect 5405 3782 5415 3834
rect 5415 3782 5461 3834
rect 5165 3780 5221 3782
rect 5245 3780 5301 3782
rect 5325 3780 5381 3782
rect 5405 3780 5461 3782
rect 5825 4378 5881 4380
rect 5905 4378 5961 4380
rect 5985 4378 6041 4380
rect 6065 4378 6121 4380
rect 5825 4326 5871 4378
rect 5871 4326 5881 4378
rect 5905 4326 5935 4378
rect 5935 4326 5947 4378
rect 5947 4326 5961 4378
rect 5985 4326 5999 4378
rect 5999 4326 6011 4378
rect 6011 4326 6041 4378
rect 6065 4326 6075 4378
rect 6075 4326 6121 4378
rect 5825 4324 5881 4326
rect 5905 4324 5961 4326
rect 5985 4324 6041 4326
rect 6065 4324 6121 4326
rect 10777 12538 10833 12540
rect 10857 12538 10913 12540
rect 10937 12538 10993 12540
rect 11017 12538 11073 12540
rect 10777 12486 10823 12538
rect 10823 12486 10833 12538
rect 10857 12486 10887 12538
rect 10887 12486 10899 12538
rect 10899 12486 10913 12538
rect 10937 12486 10951 12538
rect 10951 12486 10963 12538
rect 10963 12486 10993 12538
rect 11017 12486 11027 12538
rect 11027 12486 11073 12538
rect 10777 12484 10833 12486
rect 10857 12484 10913 12486
rect 10937 12484 10993 12486
rect 11017 12484 11073 12486
rect 8631 11994 8687 11996
rect 8711 11994 8767 11996
rect 8791 11994 8847 11996
rect 8871 11994 8927 11996
rect 8631 11942 8677 11994
rect 8677 11942 8687 11994
rect 8711 11942 8741 11994
rect 8741 11942 8753 11994
rect 8753 11942 8767 11994
rect 8791 11942 8805 11994
rect 8805 11942 8817 11994
rect 8817 11942 8847 11994
rect 8871 11942 8881 11994
rect 8881 11942 8927 11994
rect 8631 11940 8687 11942
rect 8711 11940 8767 11942
rect 8791 11940 8847 11942
rect 8871 11940 8927 11942
rect 8631 10906 8687 10908
rect 8711 10906 8767 10908
rect 8791 10906 8847 10908
rect 8871 10906 8927 10908
rect 8631 10854 8677 10906
rect 8677 10854 8687 10906
rect 8711 10854 8741 10906
rect 8741 10854 8753 10906
rect 8753 10854 8767 10906
rect 8791 10854 8805 10906
rect 8805 10854 8817 10906
rect 8817 10854 8847 10906
rect 8871 10854 8881 10906
rect 8881 10854 8927 10906
rect 8631 10852 8687 10854
rect 8711 10852 8767 10854
rect 8791 10852 8847 10854
rect 8871 10852 8927 10854
rect 8631 9818 8687 9820
rect 8711 9818 8767 9820
rect 8791 9818 8847 9820
rect 8871 9818 8927 9820
rect 8631 9766 8677 9818
rect 8677 9766 8687 9818
rect 8711 9766 8741 9818
rect 8741 9766 8753 9818
rect 8753 9766 8767 9818
rect 8791 9766 8805 9818
rect 8805 9766 8817 9818
rect 8817 9766 8847 9818
rect 8871 9766 8881 9818
rect 8881 9766 8927 9818
rect 8631 9764 8687 9766
rect 8711 9764 8767 9766
rect 8791 9764 8847 9766
rect 8871 9764 8927 9766
rect 8631 8730 8687 8732
rect 8711 8730 8767 8732
rect 8791 8730 8847 8732
rect 8871 8730 8927 8732
rect 8631 8678 8677 8730
rect 8677 8678 8687 8730
rect 8711 8678 8741 8730
rect 8741 8678 8753 8730
rect 8753 8678 8767 8730
rect 8791 8678 8805 8730
rect 8805 8678 8817 8730
rect 8817 8678 8847 8730
rect 8871 8678 8881 8730
rect 8881 8678 8927 8730
rect 8631 8676 8687 8678
rect 8711 8676 8767 8678
rect 8791 8676 8847 8678
rect 8871 8676 8927 8678
rect 7971 8186 8027 8188
rect 8051 8186 8107 8188
rect 8131 8186 8187 8188
rect 8211 8186 8267 8188
rect 7971 8134 8017 8186
rect 8017 8134 8027 8186
rect 8051 8134 8081 8186
rect 8081 8134 8093 8186
rect 8093 8134 8107 8186
rect 8131 8134 8145 8186
rect 8145 8134 8157 8186
rect 8157 8134 8187 8186
rect 8211 8134 8221 8186
rect 8221 8134 8267 8186
rect 7971 8132 8027 8134
rect 8051 8132 8107 8134
rect 8131 8132 8187 8134
rect 8211 8132 8267 8134
rect 8631 7642 8687 7644
rect 8711 7642 8767 7644
rect 8791 7642 8847 7644
rect 8871 7642 8927 7644
rect 8631 7590 8677 7642
rect 8677 7590 8687 7642
rect 8711 7590 8741 7642
rect 8741 7590 8753 7642
rect 8753 7590 8767 7642
rect 8791 7590 8805 7642
rect 8805 7590 8817 7642
rect 8817 7590 8847 7642
rect 8871 7590 8881 7642
rect 8881 7590 8927 7642
rect 8631 7588 8687 7590
rect 8711 7588 8767 7590
rect 8791 7588 8847 7590
rect 8871 7588 8927 7590
rect 7971 7098 8027 7100
rect 8051 7098 8107 7100
rect 8131 7098 8187 7100
rect 8211 7098 8267 7100
rect 7971 7046 8017 7098
rect 8017 7046 8027 7098
rect 8051 7046 8081 7098
rect 8081 7046 8093 7098
rect 8093 7046 8107 7098
rect 8131 7046 8145 7098
rect 8145 7046 8157 7098
rect 8157 7046 8187 7098
rect 8211 7046 8221 7098
rect 8221 7046 8267 7098
rect 7971 7044 8027 7046
rect 8051 7044 8107 7046
rect 8131 7044 8187 7046
rect 8211 7044 8267 7046
rect 2359 2746 2415 2748
rect 2439 2746 2495 2748
rect 2519 2746 2575 2748
rect 2599 2746 2655 2748
rect 2359 2694 2405 2746
rect 2405 2694 2415 2746
rect 2439 2694 2469 2746
rect 2469 2694 2481 2746
rect 2481 2694 2495 2746
rect 2519 2694 2533 2746
rect 2533 2694 2545 2746
rect 2545 2694 2575 2746
rect 2599 2694 2609 2746
rect 2609 2694 2655 2746
rect 2359 2692 2415 2694
rect 2439 2692 2495 2694
rect 2519 2692 2575 2694
rect 2599 2692 2655 2694
rect 5165 2746 5221 2748
rect 5245 2746 5301 2748
rect 5325 2746 5381 2748
rect 5405 2746 5461 2748
rect 5165 2694 5211 2746
rect 5211 2694 5221 2746
rect 5245 2694 5275 2746
rect 5275 2694 5287 2746
rect 5287 2694 5301 2746
rect 5325 2694 5339 2746
rect 5339 2694 5351 2746
rect 5351 2694 5381 2746
rect 5405 2694 5415 2746
rect 5415 2694 5461 2746
rect 5165 2692 5221 2694
rect 5245 2692 5301 2694
rect 5325 2692 5381 2694
rect 5405 2692 5461 2694
rect 5825 3290 5881 3292
rect 5905 3290 5961 3292
rect 5985 3290 6041 3292
rect 6065 3290 6121 3292
rect 5825 3238 5871 3290
rect 5871 3238 5881 3290
rect 5905 3238 5935 3290
rect 5935 3238 5947 3290
rect 5947 3238 5961 3290
rect 5985 3238 5999 3290
rect 5999 3238 6011 3290
rect 6011 3238 6041 3290
rect 6065 3238 6075 3290
rect 6075 3238 6121 3290
rect 5825 3236 5881 3238
rect 5905 3236 5961 3238
rect 5985 3236 6041 3238
rect 6065 3236 6121 3238
rect 7971 6010 8027 6012
rect 8051 6010 8107 6012
rect 8131 6010 8187 6012
rect 8211 6010 8267 6012
rect 7971 5958 8017 6010
rect 8017 5958 8027 6010
rect 8051 5958 8081 6010
rect 8081 5958 8093 6010
rect 8093 5958 8107 6010
rect 8131 5958 8145 6010
rect 8145 5958 8157 6010
rect 8157 5958 8187 6010
rect 8211 5958 8221 6010
rect 8221 5958 8267 6010
rect 7971 5956 8027 5958
rect 8051 5956 8107 5958
rect 8131 5956 8187 5958
rect 8211 5956 8267 5958
rect 8631 6554 8687 6556
rect 8711 6554 8767 6556
rect 8791 6554 8847 6556
rect 8871 6554 8927 6556
rect 8631 6502 8677 6554
rect 8677 6502 8687 6554
rect 8711 6502 8741 6554
rect 8741 6502 8753 6554
rect 8753 6502 8767 6554
rect 8791 6502 8805 6554
rect 8805 6502 8817 6554
rect 8817 6502 8847 6554
rect 8871 6502 8881 6554
rect 8881 6502 8927 6554
rect 8631 6500 8687 6502
rect 8711 6500 8767 6502
rect 8791 6500 8847 6502
rect 8871 6500 8927 6502
rect 7971 4922 8027 4924
rect 8051 4922 8107 4924
rect 8131 4922 8187 4924
rect 8211 4922 8267 4924
rect 7971 4870 8017 4922
rect 8017 4870 8027 4922
rect 8051 4870 8081 4922
rect 8081 4870 8093 4922
rect 8093 4870 8107 4922
rect 8131 4870 8145 4922
rect 8145 4870 8157 4922
rect 8157 4870 8187 4922
rect 8211 4870 8221 4922
rect 8221 4870 8267 4922
rect 7971 4868 8027 4870
rect 8051 4868 8107 4870
rect 8131 4868 8187 4870
rect 8211 4868 8267 4870
rect 8631 5466 8687 5468
rect 8711 5466 8767 5468
rect 8791 5466 8847 5468
rect 8871 5466 8927 5468
rect 8631 5414 8677 5466
rect 8677 5414 8687 5466
rect 8711 5414 8741 5466
rect 8741 5414 8753 5466
rect 8753 5414 8767 5466
rect 8791 5414 8805 5466
rect 8805 5414 8817 5466
rect 8817 5414 8847 5466
rect 8871 5414 8881 5466
rect 8881 5414 8927 5466
rect 8631 5412 8687 5414
rect 8711 5412 8767 5414
rect 8791 5412 8847 5414
rect 8871 5412 8927 5414
rect 10777 11450 10833 11452
rect 10857 11450 10913 11452
rect 10937 11450 10993 11452
rect 11017 11450 11073 11452
rect 10777 11398 10823 11450
rect 10823 11398 10833 11450
rect 10857 11398 10887 11450
rect 10887 11398 10899 11450
rect 10899 11398 10913 11450
rect 10937 11398 10951 11450
rect 10951 11398 10963 11450
rect 10963 11398 10993 11450
rect 11017 11398 11027 11450
rect 11027 11398 11073 11450
rect 10777 11396 10833 11398
rect 10857 11396 10913 11398
rect 10937 11396 10993 11398
rect 11017 11396 11073 11398
rect 11437 11994 11493 11996
rect 11517 11994 11573 11996
rect 11597 11994 11653 11996
rect 11677 11994 11733 11996
rect 11437 11942 11483 11994
rect 11483 11942 11493 11994
rect 11517 11942 11547 11994
rect 11547 11942 11559 11994
rect 11559 11942 11573 11994
rect 11597 11942 11611 11994
rect 11611 11942 11623 11994
rect 11623 11942 11653 11994
rect 11677 11942 11687 11994
rect 11687 11942 11733 11994
rect 11437 11940 11493 11942
rect 11517 11940 11573 11942
rect 11597 11940 11653 11942
rect 11677 11940 11733 11942
rect 11437 10906 11493 10908
rect 11517 10906 11573 10908
rect 11597 10906 11653 10908
rect 11677 10906 11733 10908
rect 11437 10854 11483 10906
rect 11483 10854 11493 10906
rect 11517 10854 11547 10906
rect 11547 10854 11559 10906
rect 11559 10854 11573 10906
rect 11597 10854 11611 10906
rect 11611 10854 11623 10906
rect 11623 10854 11653 10906
rect 11677 10854 11687 10906
rect 11687 10854 11733 10906
rect 11437 10852 11493 10854
rect 11517 10852 11573 10854
rect 11597 10852 11653 10854
rect 11677 10852 11733 10854
rect 10777 10362 10833 10364
rect 10857 10362 10913 10364
rect 10937 10362 10993 10364
rect 11017 10362 11073 10364
rect 10777 10310 10823 10362
rect 10823 10310 10833 10362
rect 10857 10310 10887 10362
rect 10887 10310 10899 10362
rect 10899 10310 10913 10362
rect 10937 10310 10951 10362
rect 10951 10310 10963 10362
rect 10963 10310 10993 10362
rect 11017 10310 11027 10362
rect 11027 10310 11073 10362
rect 10777 10308 10833 10310
rect 10857 10308 10913 10310
rect 10937 10308 10993 10310
rect 11017 10308 11073 10310
rect 10777 9274 10833 9276
rect 10857 9274 10913 9276
rect 10937 9274 10993 9276
rect 11017 9274 11073 9276
rect 10777 9222 10823 9274
rect 10823 9222 10833 9274
rect 10857 9222 10887 9274
rect 10887 9222 10899 9274
rect 10899 9222 10913 9274
rect 10937 9222 10951 9274
rect 10951 9222 10963 9274
rect 10963 9222 10993 9274
rect 11017 9222 11027 9274
rect 11027 9222 11073 9274
rect 10777 9220 10833 9222
rect 10857 9220 10913 9222
rect 10937 9220 10993 9222
rect 11017 9220 11073 9222
rect 11437 9818 11493 9820
rect 11517 9818 11573 9820
rect 11597 9818 11653 9820
rect 11677 9818 11733 9820
rect 11437 9766 11483 9818
rect 11483 9766 11493 9818
rect 11517 9766 11547 9818
rect 11547 9766 11559 9818
rect 11559 9766 11573 9818
rect 11597 9766 11611 9818
rect 11611 9766 11623 9818
rect 11623 9766 11653 9818
rect 11677 9766 11687 9818
rect 11687 9766 11733 9818
rect 11437 9764 11493 9766
rect 11517 9764 11573 9766
rect 11597 9764 11653 9766
rect 11677 9764 11733 9766
rect 11978 9560 12034 9616
rect 10777 8186 10833 8188
rect 10857 8186 10913 8188
rect 10937 8186 10993 8188
rect 11017 8186 11073 8188
rect 10777 8134 10823 8186
rect 10823 8134 10833 8186
rect 10857 8134 10887 8186
rect 10887 8134 10899 8186
rect 10899 8134 10913 8186
rect 10937 8134 10951 8186
rect 10951 8134 10963 8186
rect 10963 8134 10993 8186
rect 11017 8134 11027 8186
rect 11027 8134 11073 8186
rect 10777 8132 10833 8134
rect 10857 8132 10913 8134
rect 10937 8132 10993 8134
rect 11017 8132 11073 8134
rect 10777 7098 10833 7100
rect 10857 7098 10913 7100
rect 10937 7098 10993 7100
rect 11017 7098 11073 7100
rect 10777 7046 10823 7098
rect 10823 7046 10833 7098
rect 10857 7046 10887 7098
rect 10887 7046 10899 7098
rect 10899 7046 10913 7098
rect 10937 7046 10951 7098
rect 10951 7046 10963 7098
rect 10963 7046 10993 7098
rect 11017 7046 11027 7098
rect 11027 7046 11073 7098
rect 10777 7044 10833 7046
rect 10857 7044 10913 7046
rect 10937 7044 10993 7046
rect 11017 7044 11073 7046
rect 8631 4378 8687 4380
rect 8711 4378 8767 4380
rect 8791 4378 8847 4380
rect 8871 4378 8927 4380
rect 8631 4326 8677 4378
rect 8677 4326 8687 4378
rect 8711 4326 8741 4378
rect 8741 4326 8753 4378
rect 8753 4326 8767 4378
rect 8791 4326 8805 4378
rect 8805 4326 8817 4378
rect 8817 4326 8847 4378
rect 8871 4326 8881 4378
rect 8881 4326 8927 4378
rect 8631 4324 8687 4326
rect 8711 4324 8767 4326
rect 8791 4324 8847 4326
rect 8871 4324 8927 4326
rect 7971 3834 8027 3836
rect 8051 3834 8107 3836
rect 8131 3834 8187 3836
rect 8211 3834 8267 3836
rect 7971 3782 8017 3834
rect 8017 3782 8027 3834
rect 8051 3782 8081 3834
rect 8081 3782 8093 3834
rect 8093 3782 8107 3834
rect 8131 3782 8145 3834
rect 8145 3782 8157 3834
rect 8157 3782 8187 3834
rect 8211 3782 8221 3834
rect 8221 3782 8267 3834
rect 7971 3780 8027 3782
rect 8051 3780 8107 3782
rect 8131 3780 8187 3782
rect 8211 3780 8267 3782
rect 8631 3290 8687 3292
rect 8711 3290 8767 3292
rect 8791 3290 8847 3292
rect 8871 3290 8927 3292
rect 8631 3238 8677 3290
rect 8677 3238 8687 3290
rect 8711 3238 8741 3290
rect 8741 3238 8753 3290
rect 8753 3238 8767 3290
rect 8791 3238 8805 3290
rect 8805 3238 8817 3290
rect 8817 3238 8847 3290
rect 8871 3238 8881 3290
rect 8881 3238 8927 3290
rect 8631 3236 8687 3238
rect 8711 3236 8767 3238
rect 8791 3236 8847 3238
rect 8871 3236 8927 3238
rect 11886 8880 11942 8936
rect 11437 8730 11493 8732
rect 11517 8730 11573 8732
rect 11597 8730 11653 8732
rect 11677 8730 11733 8732
rect 11437 8678 11483 8730
rect 11483 8678 11493 8730
rect 11517 8678 11547 8730
rect 11547 8678 11559 8730
rect 11559 8678 11573 8730
rect 11597 8678 11611 8730
rect 11611 8678 11623 8730
rect 11623 8678 11653 8730
rect 11677 8678 11687 8730
rect 11687 8678 11733 8730
rect 11437 8676 11493 8678
rect 11517 8676 11573 8678
rect 11597 8676 11653 8678
rect 11677 8676 11733 8678
rect 11437 7642 11493 7644
rect 11517 7642 11573 7644
rect 11597 7642 11653 7644
rect 11677 7642 11733 7644
rect 11437 7590 11483 7642
rect 11483 7590 11493 7642
rect 11517 7590 11547 7642
rect 11547 7590 11559 7642
rect 11559 7590 11573 7642
rect 11597 7590 11611 7642
rect 11611 7590 11623 7642
rect 11623 7590 11653 7642
rect 11677 7590 11687 7642
rect 11687 7590 11733 7642
rect 11437 7588 11493 7590
rect 11517 7588 11573 7590
rect 11597 7588 11653 7590
rect 11677 7588 11733 7590
rect 11437 6554 11493 6556
rect 11517 6554 11573 6556
rect 11597 6554 11653 6556
rect 11677 6554 11733 6556
rect 11437 6502 11483 6554
rect 11483 6502 11493 6554
rect 11517 6502 11547 6554
rect 11547 6502 11559 6554
rect 11559 6502 11573 6554
rect 11597 6502 11611 6554
rect 11611 6502 11623 6554
rect 11623 6502 11653 6554
rect 11677 6502 11687 6554
rect 11687 6502 11733 6554
rect 11437 6500 11493 6502
rect 11517 6500 11573 6502
rect 11597 6500 11653 6502
rect 11677 6500 11733 6502
rect 10777 6010 10833 6012
rect 10857 6010 10913 6012
rect 10937 6010 10993 6012
rect 11017 6010 11073 6012
rect 10777 5958 10823 6010
rect 10823 5958 10833 6010
rect 10857 5958 10887 6010
rect 10887 5958 10899 6010
rect 10899 5958 10913 6010
rect 10937 5958 10951 6010
rect 10951 5958 10963 6010
rect 10963 5958 10993 6010
rect 11017 5958 11027 6010
rect 11027 5958 11073 6010
rect 10777 5956 10833 5958
rect 10857 5956 10913 5958
rect 10937 5956 10993 5958
rect 11017 5956 11073 5958
rect 11886 6180 11942 6216
rect 11886 6160 11888 6180
rect 11888 6160 11940 6180
rect 11940 6160 11942 6180
rect 11978 5480 12034 5536
rect 11437 5466 11493 5468
rect 11517 5466 11573 5468
rect 11597 5466 11653 5468
rect 11677 5466 11733 5468
rect 11437 5414 11483 5466
rect 11483 5414 11493 5466
rect 11517 5414 11547 5466
rect 11547 5414 11559 5466
rect 11559 5414 11573 5466
rect 11597 5414 11611 5466
rect 11611 5414 11623 5466
rect 11623 5414 11653 5466
rect 11677 5414 11687 5466
rect 11687 5414 11733 5466
rect 11437 5412 11493 5414
rect 11517 5412 11573 5414
rect 11597 5412 11653 5414
rect 11677 5412 11733 5414
rect 10777 4922 10833 4924
rect 10857 4922 10913 4924
rect 10937 4922 10993 4924
rect 11017 4922 11073 4924
rect 10777 4870 10823 4922
rect 10823 4870 10833 4922
rect 10857 4870 10887 4922
rect 10887 4870 10899 4922
rect 10899 4870 10913 4922
rect 10937 4870 10951 4922
rect 10951 4870 10963 4922
rect 10963 4870 10993 4922
rect 11017 4870 11027 4922
rect 11027 4870 11073 4922
rect 10777 4868 10833 4870
rect 10857 4868 10913 4870
rect 10937 4868 10993 4870
rect 11017 4868 11073 4870
rect 11978 4800 12034 4856
rect 11437 4378 11493 4380
rect 11517 4378 11573 4380
rect 11597 4378 11653 4380
rect 11677 4378 11733 4380
rect 11437 4326 11483 4378
rect 11483 4326 11493 4378
rect 11517 4326 11547 4378
rect 11547 4326 11559 4378
rect 11559 4326 11573 4378
rect 11597 4326 11611 4378
rect 11611 4326 11623 4378
rect 11623 4326 11653 4378
rect 11677 4326 11687 4378
rect 11687 4326 11733 4378
rect 11437 4324 11493 4326
rect 11517 4324 11573 4326
rect 11597 4324 11653 4326
rect 11677 4324 11733 4326
rect 10777 3834 10833 3836
rect 10857 3834 10913 3836
rect 10937 3834 10993 3836
rect 11017 3834 11073 3836
rect 10777 3782 10823 3834
rect 10823 3782 10833 3834
rect 10857 3782 10887 3834
rect 10887 3782 10899 3834
rect 10899 3782 10913 3834
rect 10937 3782 10951 3834
rect 10951 3782 10963 3834
rect 10963 3782 10993 3834
rect 11017 3782 11027 3834
rect 11027 3782 11073 3834
rect 10777 3780 10833 3782
rect 10857 3780 10913 3782
rect 10937 3780 10993 3782
rect 11017 3780 11073 3782
rect 11886 3460 11942 3496
rect 11886 3440 11888 3460
rect 11888 3440 11940 3460
rect 11940 3440 11942 3460
rect 11437 3290 11493 3292
rect 11517 3290 11573 3292
rect 11597 3290 11653 3292
rect 11677 3290 11733 3292
rect 11437 3238 11483 3290
rect 11483 3238 11493 3290
rect 11517 3238 11547 3290
rect 11547 3238 11559 3290
rect 11559 3238 11573 3290
rect 11597 3238 11611 3290
rect 11611 3238 11623 3290
rect 11623 3238 11653 3290
rect 11677 3238 11687 3290
rect 11687 3238 11733 3290
rect 11437 3236 11493 3238
rect 11517 3236 11573 3238
rect 11597 3236 11653 3238
rect 11677 3236 11733 3238
rect 7971 2746 8027 2748
rect 8051 2746 8107 2748
rect 8131 2746 8187 2748
rect 8211 2746 8267 2748
rect 7971 2694 8017 2746
rect 8017 2694 8027 2746
rect 8051 2694 8081 2746
rect 8081 2694 8093 2746
rect 8093 2694 8107 2746
rect 8131 2694 8145 2746
rect 8145 2694 8157 2746
rect 8157 2694 8187 2746
rect 8211 2694 8221 2746
rect 8221 2694 8267 2746
rect 7971 2692 8027 2694
rect 8051 2692 8107 2694
rect 8131 2692 8187 2694
rect 8211 2692 8267 2694
rect 10777 2746 10833 2748
rect 10857 2746 10913 2748
rect 10937 2746 10993 2748
rect 11017 2746 11073 2748
rect 10777 2694 10823 2746
rect 10823 2694 10833 2746
rect 10857 2694 10887 2746
rect 10887 2694 10899 2746
rect 10899 2694 10913 2746
rect 10937 2694 10951 2746
rect 10951 2694 10963 2746
rect 10963 2694 10993 2746
rect 11017 2694 11027 2746
rect 11027 2694 11073 2746
rect 10777 2692 10833 2694
rect 10857 2692 10913 2694
rect 10937 2692 10993 2694
rect 11017 2692 11073 2694
rect 3019 2202 3075 2204
rect 3099 2202 3155 2204
rect 3179 2202 3235 2204
rect 3259 2202 3315 2204
rect 3019 2150 3065 2202
rect 3065 2150 3075 2202
rect 3099 2150 3129 2202
rect 3129 2150 3141 2202
rect 3141 2150 3155 2202
rect 3179 2150 3193 2202
rect 3193 2150 3205 2202
rect 3205 2150 3235 2202
rect 3259 2150 3269 2202
rect 3269 2150 3315 2202
rect 3019 2148 3075 2150
rect 3099 2148 3155 2150
rect 3179 2148 3235 2150
rect 3259 2148 3315 2150
rect 5825 2202 5881 2204
rect 5905 2202 5961 2204
rect 5985 2202 6041 2204
rect 6065 2202 6121 2204
rect 5825 2150 5871 2202
rect 5871 2150 5881 2202
rect 5905 2150 5935 2202
rect 5935 2150 5947 2202
rect 5947 2150 5961 2202
rect 5985 2150 5999 2202
rect 5999 2150 6011 2202
rect 6011 2150 6041 2202
rect 6065 2150 6075 2202
rect 6075 2150 6121 2202
rect 5825 2148 5881 2150
rect 5905 2148 5961 2150
rect 5985 2148 6041 2150
rect 6065 2148 6121 2150
rect 8631 2202 8687 2204
rect 8711 2202 8767 2204
rect 8791 2202 8847 2204
rect 8871 2202 8927 2204
rect 8631 2150 8677 2202
rect 8677 2150 8687 2202
rect 8711 2150 8741 2202
rect 8741 2150 8753 2202
rect 8753 2150 8767 2202
rect 8791 2150 8805 2202
rect 8805 2150 8817 2202
rect 8817 2150 8847 2202
rect 8871 2150 8881 2202
rect 8881 2150 8927 2202
rect 8631 2148 8687 2150
rect 8711 2148 8767 2150
rect 8791 2148 8847 2150
rect 8871 2148 8927 2150
rect 11437 2202 11493 2204
rect 11517 2202 11573 2204
rect 11597 2202 11653 2204
rect 11677 2202 11733 2204
rect 11437 2150 11483 2202
rect 11483 2150 11493 2202
rect 11517 2150 11547 2202
rect 11547 2150 11559 2202
rect 11559 2150 11573 2202
rect 11597 2150 11611 2202
rect 11611 2150 11623 2202
rect 11623 2150 11653 2202
rect 11677 2150 11687 2202
rect 11687 2150 11733 2202
rect 11437 2148 11493 2150
rect 11517 2148 11573 2150
rect 11597 2148 11653 2150
rect 11677 2148 11733 2150
<< metal3 >>
rect 3009 13088 3325 13089
rect 3009 13024 3015 13088
rect 3079 13024 3095 13088
rect 3159 13024 3175 13088
rect 3239 13024 3255 13088
rect 3319 13024 3325 13088
rect 3009 13023 3325 13024
rect 5815 13088 6131 13089
rect 5815 13024 5821 13088
rect 5885 13024 5901 13088
rect 5965 13024 5981 13088
rect 6045 13024 6061 13088
rect 6125 13024 6131 13088
rect 5815 13023 6131 13024
rect 8621 13088 8937 13089
rect 8621 13024 8627 13088
rect 8691 13024 8707 13088
rect 8771 13024 8787 13088
rect 8851 13024 8867 13088
rect 8931 13024 8937 13088
rect 8621 13023 8937 13024
rect 11427 13088 11743 13089
rect 11427 13024 11433 13088
rect 11497 13024 11513 13088
rect 11577 13024 11593 13088
rect 11657 13024 11673 13088
rect 11737 13024 11743 13088
rect 11427 13023 11743 13024
rect 2349 12544 2665 12545
rect 2349 12480 2355 12544
rect 2419 12480 2435 12544
rect 2499 12480 2515 12544
rect 2579 12480 2595 12544
rect 2659 12480 2665 12544
rect 2349 12479 2665 12480
rect 5155 12544 5471 12545
rect 5155 12480 5161 12544
rect 5225 12480 5241 12544
rect 5305 12480 5321 12544
rect 5385 12480 5401 12544
rect 5465 12480 5471 12544
rect 5155 12479 5471 12480
rect 7961 12544 8277 12545
rect 7961 12480 7967 12544
rect 8031 12480 8047 12544
rect 8111 12480 8127 12544
rect 8191 12480 8207 12544
rect 8271 12480 8277 12544
rect 7961 12479 8277 12480
rect 10767 12544 11083 12545
rect 10767 12480 10773 12544
rect 10837 12480 10853 12544
rect 10917 12480 10933 12544
rect 10997 12480 11013 12544
rect 11077 12480 11083 12544
rect 10767 12479 11083 12480
rect 3009 12000 3325 12001
rect 3009 11936 3015 12000
rect 3079 11936 3095 12000
rect 3159 11936 3175 12000
rect 3239 11936 3255 12000
rect 3319 11936 3325 12000
rect 3009 11935 3325 11936
rect 5815 12000 6131 12001
rect 5815 11936 5821 12000
rect 5885 11936 5901 12000
rect 5965 11936 5981 12000
rect 6045 11936 6061 12000
rect 6125 11936 6131 12000
rect 5815 11935 6131 11936
rect 8621 12000 8937 12001
rect 8621 11936 8627 12000
rect 8691 11936 8707 12000
rect 8771 11936 8787 12000
rect 8851 11936 8867 12000
rect 8931 11936 8937 12000
rect 8621 11935 8937 11936
rect 11427 12000 11743 12001
rect 11427 11936 11433 12000
rect 11497 11936 11513 12000
rect 11577 11936 11593 12000
rect 11657 11936 11673 12000
rect 11737 11936 11743 12000
rect 11427 11935 11743 11936
rect 0 11658 800 11688
rect 4102 11658 4108 11660
rect 0 11598 4108 11658
rect 0 11568 800 11598
rect 4102 11596 4108 11598
rect 4172 11596 4178 11660
rect 2349 11456 2665 11457
rect 2349 11392 2355 11456
rect 2419 11392 2435 11456
rect 2499 11392 2515 11456
rect 2579 11392 2595 11456
rect 2659 11392 2665 11456
rect 2349 11391 2665 11392
rect 5155 11456 5471 11457
rect 5155 11392 5161 11456
rect 5225 11392 5241 11456
rect 5305 11392 5321 11456
rect 5385 11392 5401 11456
rect 5465 11392 5471 11456
rect 5155 11391 5471 11392
rect 7961 11456 8277 11457
rect 7961 11392 7967 11456
rect 8031 11392 8047 11456
rect 8111 11392 8127 11456
rect 8191 11392 8207 11456
rect 8271 11392 8277 11456
rect 7961 11391 8277 11392
rect 10767 11456 11083 11457
rect 10767 11392 10773 11456
rect 10837 11392 10853 11456
rect 10917 11392 10933 11456
rect 10997 11392 11013 11456
rect 11077 11392 11083 11456
rect 10767 11391 11083 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 3009 10912 3325 10913
rect 3009 10848 3015 10912
rect 3079 10848 3095 10912
rect 3159 10848 3175 10912
rect 3239 10848 3255 10912
rect 3319 10848 3325 10912
rect 3009 10847 3325 10848
rect 5815 10912 6131 10913
rect 5815 10848 5821 10912
rect 5885 10848 5901 10912
rect 5965 10848 5981 10912
rect 6045 10848 6061 10912
rect 6125 10848 6131 10912
rect 5815 10847 6131 10848
rect 8621 10912 8937 10913
rect 8621 10848 8627 10912
rect 8691 10848 8707 10912
rect 8771 10848 8787 10912
rect 8851 10848 8867 10912
rect 8931 10848 8937 10912
rect 8621 10847 8937 10848
rect 11427 10912 11743 10913
rect 11427 10848 11433 10912
rect 11497 10848 11513 10912
rect 11577 10848 11593 10912
rect 11657 10848 11673 10912
rect 11737 10848 11743 10912
rect 11427 10847 11743 10848
rect 2349 10368 2665 10369
rect 0 10298 800 10328
rect 2349 10304 2355 10368
rect 2419 10304 2435 10368
rect 2499 10304 2515 10368
rect 2579 10304 2595 10368
rect 2659 10304 2665 10368
rect 2349 10303 2665 10304
rect 5155 10368 5471 10369
rect 5155 10304 5161 10368
rect 5225 10304 5241 10368
rect 5305 10304 5321 10368
rect 5385 10304 5401 10368
rect 5465 10304 5471 10368
rect 5155 10303 5471 10304
rect 7961 10368 8277 10369
rect 7961 10304 7967 10368
rect 8031 10304 8047 10368
rect 8111 10304 8127 10368
rect 8191 10304 8207 10368
rect 8271 10304 8277 10368
rect 7961 10303 8277 10304
rect 10767 10368 11083 10369
rect 10767 10304 10773 10368
rect 10837 10304 10853 10368
rect 10917 10304 10933 10368
rect 10997 10304 11013 10368
rect 11077 10304 11083 10368
rect 10767 10303 11083 10304
rect 1301 10298 1367 10301
rect 0 10296 1367 10298
rect 0 10240 1306 10296
rect 1362 10240 1367 10296
rect 0 10238 1367 10240
rect 0 10208 800 10238
rect 1301 10235 1367 10238
rect 3009 9824 3325 9825
rect 3009 9760 3015 9824
rect 3079 9760 3095 9824
rect 3159 9760 3175 9824
rect 3239 9760 3255 9824
rect 3319 9760 3325 9824
rect 3009 9759 3325 9760
rect 5815 9824 6131 9825
rect 5815 9760 5821 9824
rect 5885 9760 5901 9824
rect 5965 9760 5981 9824
rect 6045 9760 6061 9824
rect 6125 9760 6131 9824
rect 5815 9759 6131 9760
rect 8621 9824 8937 9825
rect 8621 9760 8627 9824
rect 8691 9760 8707 9824
rect 8771 9760 8787 9824
rect 8851 9760 8867 9824
rect 8931 9760 8937 9824
rect 8621 9759 8937 9760
rect 11427 9824 11743 9825
rect 11427 9760 11433 9824
rect 11497 9760 11513 9824
rect 11577 9760 11593 9824
rect 11657 9760 11673 9824
rect 11737 9760 11743 9824
rect 11427 9759 11743 9760
rect 11973 9618 12039 9621
rect 12699 9618 13499 9648
rect 11973 9616 13499 9618
rect 11973 9560 11978 9616
rect 12034 9560 13499 9616
rect 11973 9558 13499 9560
rect 11973 9555 12039 9558
rect 12699 9528 13499 9558
rect 2349 9280 2665 9281
rect 2349 9216 2355 9280
rect 2419 9216 2435 9280
rect 2499 9216 2515 9280
rect 2579 9216 2595 9280
rect 2659 9216 2665 9280
rect 2349 9215 2665 9216
rect 5155 9280 5471 9281
rect 5155 9216 5161 9280
rect 5225 9216 5241 9280
rect 5305 9216 5321 9280
rect 5385 9216 5401 9280
rect 5465 9216 5471 9280
rect 5155 9215 5471 9216
rect 7961 9280 8277 9281
rect 7961 9216 7967 9280
rect 8031 9216 8047 9280
rect 8111 9216 8127 9280
rect 8191 9216 8207 9280
rect 8271 9216 8277 9280
rect 7961 9215 8277 9216
rect 10767 9280 11083 9281
rect 10767 9216 10773 9280
rect 10837 9216 10853 9280
rect 10917 9216 10933 9280
rect 10997 9216 11013 9280
rect 11077 9216 11083 9280
rect 10767 9215 11083 9216
rect 11881 8938 11947 8941
rect 12699 8938 13499 8968
rect 11881 8936 13499 8938
rect 11881 8880 11886 8936
rect 11942 8880 13499 8936
rect 11881 8878 13499 8880
rect 11881 8875 11947 8878
rect 12699 8848 13499 8878
rect 3009 8736 3325 8737
rect 3009 8672 3015 8736
rect 3079 8672 3095 8736
rect 3159 8672 3175 8736
rect 3239 8672 3255 8736
rect 3319 8672 3325 8736
rect 3009 8671 3325 8672
rect 5815 8736 6131 8737
rect 5815 8672 5821 8736
rect 5885 8672 5901 8736
rect 5965 8672 5981 8736
rect 6045 8672 6061 8736
rect 6125 8672 6131 8736
rect 5815 8671 6131 8672
rect 8621 8736 8937 8737
rect 8621 8672 8627 8736
rect 8691 8672 8707 8736
rect 8771 8672 8787 8736
rect 8851 8672 8867 8736
rect 8931 8672 8937 8736
rect 8621 8671 8937 8672
rect 11427 8736 11743 8737
rect 11427 8672 11433 8736
rect 11497 8672 11513 8736
rect 11577 8672 11593 8736
rect 11657 8672 11673 8736
rect 11737 8672 11743 8736
rect 11427 8671 11743 8672
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 4102 8196 4108 8260
rect 4172 8258 4178 8260
rect 4245 8258 4311 8261
rect 4172 8256 4311 8258
rect 4172 8200 4250 8256
rect 4306 8200 4311 8256
rect 4172 8198 4311 8200
rect 4172 8196 4178 8198
rect 4245 8195 4311 8198
rect 2349 8192 2665 8193
rect 2349 8128 2355 8192
rect 2419 8128 2435 8192
rect 2499 8128 2515 8192
rect 2579 8128 2595 8192
rect 2659 8128 2665 8192
rect 2349 8127 2665 8128
rect 5155 8192 5471 8193
rect 5155 8128 5161 8192
rect 5225 8128 5241 8192
rect 5305 8128 5321 8192
rect 5385 8128 5401 8192
rect 5465 8128 5471 8192
rect 5155 8127 5471 8128
rect 7961 8192 8277 8193
rect 7961 8128 7967 8192
rect 8031 8128 8047 8192
rect 8111 8128 8127 8192
rect 8191 8128 8207 8192
rect 8271 8128 8277 8192
rect 7961 8127 8277 8128
rect 10767 8192 11083 8193
rect 10767 8128 10773 8192
rect 10837 8128 10853 8192
rect 10917 8128 10933 8192
rect 10997 8128 11013 8192
rect 11077 8128 11083 8192
rect 10767 8127 11083 8128
rect 3009 7648 3325 7649
rect 3009 7584 3015 7648
rect 3079 7584 3095 7648
rect 3159 7584 3175 7648
rect 3239 7584 3255 7648
rect 3319 7584 3325 7648
rect 3009 7583 3325 7584
rect 5815 7648 6131 7649
rect 5815 7584 5821 7648
rect 5885 7584 5901 7648
rect 5965 7584 5981 7648
rect 6045 7584 6061 7648
rect 6125 7584 6131 7648
rect 5815 7583 6131 7584
rect 8621 7648 8937 7649
rect 8621 7584 8627 7648
rect 8691 7584 8707 7648
rect 8771 7584 8787 7648
rect 8851 7584 8867 7648
rect 8931 7584 8937 7648
rect 8621 7583 8937 7584
rect 11427 7648 11743 7649
rect 11427 7584 11433 7648
rect 11497 7584 11513 7648
rect 11577 7584 11593 7648
rect 11657 7584 11673 7648
rect 11737 7584 11743 7648
rect 11427 7583 11743 7584
rect 2349 7104 2665 7105
rect 2349 7040 2355 7104
rect 2419 7040 2435 7104
rect 2499 7040 2515 7104
rect 2579 7040 2595 7104
rect 2659 7040 2665 7104
rect 2349 7039 2665 7040
rect 5155 7104 5471 7105
rect 5155 7040 5161 7104
rect 5225 7040 5241 7104
rect 5305 7040 5321 7104
rect 5385 7040 5401 7104
rect 5465 7040 5471 7104
rect 5155 7039 5471 7040
rect 7961 7104 8277 7105
rect 7961 7040 7967 7104
rect 8031 7040 8047 7104
rect 8111 7040 8127 7104
rect 8191 7040 8207 7104
rect 8271 7040 8277 7104
rect 7961 7039 8277 7040
rect 10767 7104 11083 7105
rect 10767 7040 10773 7104
rect 10837 7040 10853 7104
rect 10917 7040 10933 7104
rect 10997 7040 11013 7104
rect 11077 7040 11083 7104
rect 10767 7039 11083 7040
rect 3009 6560 3325 6561
rect 3009 6496 3015 6560
rect 3079 6496 3095 6560
rect 3159 6496 3175 6560
rect 3239 6496 3255 6560
rect 3319 6496 3325 6560
rect 3009 6495 3325 6496
rect 5815 6560 6131 6561
rect 5815 6496 5821 6560
rect 5885 6496 5901 6560
rect 5965 6496 5981 6560
rect 6045 6496 6061 6560
rect 6125 6496 6131 6560
rect 5815 6495 6131 6496
rect 8621 6560 8937 6561
rect 8621 6496 8627 6560
rect 8691 6496 8707 6560
rect 8771 6496 8787 6560
rect 8851 6496 8867 6560
rect 8931 6496 8937 6560
rect 8621 6495 8937 6496
rect 11427 6560 11743 6561
rect 11427 6496 11433 6560
rect 11497 6496 11513 6560
rect 11577 6496 11593 6560
rect 11657 6496 11673 6560
rect 11737 6496 11743 6560
rect 11427 6495 11743 6496
rect 11881 6218 11947 6221
rect 12699 6218 13499 6248
rect 11881 6216 13499 6218
rect 11881 6160 11886 6216
rect 11942 6160 13499 6216
rect 11881 6158 13499 6160
rect 11881 6155 11947 6158
rect 12699 6128 13499 6158
rect 2349 6016 2665 6017
rect 2349 5952 2355 6016
rect 2419 5952 2435 6016
rect 2499 5952 2515 6016
rect 2579 5952 2595 6016
rect 2659 5952 2665 6016
rect 2349 5951 2665 5952
rect 5155 6016 5471 6017
rect 5155 5952 5161 6016
rect 5225 5952 5241 6016
rect 5305 5952 5321 6016
rect 5385 5952 5401 6016
rect 5465 5952 5471 6016
rect 5155 5951 5471 5952
rect 7961 6016 8277 6017
rect 7961 5952 7967 6016
rect 8031 5952 8047 6016
rect 8111 5952 8127 6016
rect 8191 5952 8207 6016
rect 8271 5952 8277 6016
rect 7961 5951 8277 5952
rect 10767 6016 11083 6017
rect 10767 5952 10773 6016
rect 10837 5952 10853 6016
rect 10917 5952 10933 6016
rect 10997 5952 11013 6016
rect 11077 5952 11083 6016
rect 10767 5951 11083 5952
rect 11973 5538 12039 5541
rect 12699 5538 13499 5568
rect 11973 5536 13499 5538
rect 11973 5480 11978 5536
rect 12034 5480 13499 5536
rect 11973 5478 13499 5480
rect 11973 5475 12039 5478
rect 3009 5472 3325 5473
rect 3009 5408 3015 5472
rect 3079 5408 3095 5472
rect 3159 5408 3175 5472
rect 3239 5408 3255 5472
rect 3319 5408 3325 5472
rect 3009 5407 3325 5408
rect 5815 5472 6131 5473
rect 5815 5408 5821 5472
rect 5885 5408 5901 5472
rect 5965 5408 5981 5472
rect 6045 5408 6061 5472
rect 6125 5408 6131 5472
rect 5815 5407 6131 5408
rect 8621 5472 8937 5473
rect 8621 5408 8627 5472
rect 8691 5408 8707 5472
rect 8771 5408 8787 5472
rect 8851 5408 8867 5472
rect 8931 5408 8937 5472
rect 8621 5407 8937 5408
rect 11427 5472 11743 5473
rect 11427 5408 11433 5472
rect 11497 5408 11513 5472
rect 11577 5408 11593 5472
rect 11657 5408 11673 5472
rect 11737 5408 11743 5472
rect 12699 5448 13499 5478
rect 11427 5407 11743 5408
rect 2349 4928 2665 4929
rect 2349 4864 2355 4928
rect 2419 4864 2435 4928
rect 2499 4864 2515 4928
rect 2579 4864 2595 4928
rect 2659 4864 2665 4928
rect 2349 4863 2665 4864
rect 5155 4928 5471 4929
rect 5155 4864 5161 4928
rect 5225 4864 5241 4928
rect 5305 4864 5321 4928
rect 5385 4864 5401 4928
rect 5465 4864 5471 4928
rect 5155 4863 5471 4864
rect 7961 4928 8277 4929
rect 7961 4864 7967 4928
rect 8031 4864 8047 4928
rect 8111 4864 8127 4928
rect 8191 4864 8207 4928
rect 8271 4864 8277 4928
rect 7961 4863 8277 4864
rect 10767 4928 11083 4929
rect 10767 4864 10773 4928
rect 10837 4864 10853 4928
rect 10917 4864 10933 4928
rect 10997 4864 11013 4928
rect 11077 4864 11083 4928
rect 10767 4863 11083 4864
rect 11973 4858 12039 4861
rect 12699 4858 13499 4888
rect 11973 4856 13499 4858
rect 11973 4800 11978 4856
rect 12034 4800 13499 4856
rect 11973 4798 13499 4800
rect 11973 4795 12039 4798
rect 12699 4768 13499 4798
rect 3009 4384 3325 4385
rect 3009 4320 3015 4384
rect 3079 4320 3095 4384
rect 3159 4320 3175 4384
rect 3239 4320 3255 4384
rect 3319 4320 3325 4384
rect 3009 4319 3325 4320
rect 5815 4384 6131 4385
rect 5815 4320 5821 4384
rect 5885 4320 5901 4384
rect 5965 4320 5981 4384
rect 6045 4320 6061 4384
rect 6125 4320 6131 4384
rect 5815 4319 6131 4320
rect 8621 4384 8937 4385
rect 8621 4320 8627 4384
rect 8691 4320 8707 4384
rect 8771 4320 8787 4384
rect 8851 4320 8867 4384
rect 8931 4320 8937 4384
rect 8621 4319 8937 4320
rect 11427 4384 11743 4385
rect 11427 4320 11433 4384
rect 11497 4320 11513 4384
rect 11577 4320 11593 4384
rect 11657 4320 11673 4384
rect 11737 4320 11743 4384
rect 11427 4319 11743 4320
rect 2349 3840 2665 3841
rect 2349 3776 2355 3840
rect 2419 3776 2435 3840
rect 2499 3776 2515 3840
rect 2579 3776 2595 3840
rect 2659 3776 2665 3840
rect 2349 3775 2665 3776
rect 5155 3840 5471 3841
rect 5155 3776 5161 3840
rect 5225 3776 5241 3840
rect 5305 3776 5321 3840
rect 5385 3776 5401 3840
rect 5465 3776 5471 3840
rect 5155 3775 5471 3776
rect 7961 3840 8277 3841
rect 7961 3776 7967 3840
rect 8031 3776 8047 3840
rect 8111 3776 8127 3840
rect 8191 3776 8207 3840
rect 8271 3776 8277 3840
rect 7961 3775 8277 3776
rect 10767 3840 11083 3841
rect 10767 3776 10773 3840
rect 10837 3776 10853 3840
rect 10917 3776 10933 3840
rect 10997 3776 11013 3840
rect 11077 3776 11083 3840
rect 10767 3775 11083 3776
rect 11881 3498 11947 3501
rect 12699 3498 13499 3528
rect 11881 3496 13499 3498
rect 11881 3440 11886 3496
rect 11942 3440 13499 3496
rect 11881 3438 13499 3440
rect 11881 3435 11947 3438
rect 12699 3408 13499 3438
rect 3009 3296 3325 3297
rect 3009 3232 3015 3296
rect 3079 3232 3095 3296
rect 3159 3232 3175 3296
rect 3239 3232 3255 3296
rect 3319 3232 3325 3296
rect 3009 3231 3325 3232
rect 5815 3296 6131 3297
rect 5815 3232 5821 3296
rect 5885 3232 5901 3296
rect 5965 3232 5981 3296
rect 6045 3232 6061 3296
rect 6125 3232 6131 3296
rect 5815 3231 6131 3232
rect 8621 3296 8937 3297
rect 8621 3232 8627 3296
rect 8691 3232 8707 3296
rect 8771 3232 8787 3296
rect 8851 3232 8867 3296
rect 8931 3232 8937 3296
rect 8621 3231 8937 3232
rect 11427 3296 11743 3297
rect 11427 3232 11433 3296
rect 11497 3232 11513 3296
rect 11577 3232 11593 3296
rect 11657 3232 11673 3296
rect 11737 3232 11743 3296
rect 11427 3231 11743 3232
rect 2349 2752 2665 2753
rect 2349 2688 2355 2752
rect 2419 2688 2435 2752
rect 2499 2688 2515 2752
rect 2579 2688 2595 2752
rect 2659 2688 2665 2752
rect 2349 2687 2665 2688
rect 5155 2752 5471 2753
rect 5155 2688 5161 2752
rect 5225 2688 5241 2752
rect 5305 2688 5321 2752
rect 5385 2688 5401 2752
rect 5465 2688 5471 2752
rect 5155 2687 5471 2688
rect 7961 2752 8277 2753
rect 7961 2688 7967 2752
rect 8031 2688 8047 2752
rect 8111 2688 8127 2752
rect 8191 2688 8207 2752
rect 8271 2688 8277 2752
rect 7961 2687 8277 2688
rect 10767 2752 11083 2753
rect 10767 2688 10773 2752
rect 10837 2688 10853 2752
rect 10917 2688 10933 2752
rect 10997 2688 11013 2752
rect 11077 2688 11083 2752
rect 10767 2687 11083 2688
rect 3009 2208 3325 2209
rect 3009 2144 3015 2208
rect 3079 2144 3095 2208
rect 3159 2144 3175 2208
rect 3239 2144 3255 2208
rect 3319 2144 3325 2208
rect 3009 2143 3325 2144
rect 5815 2208 6131 2209
rect 5815 2144 5821 2208
rect 5885 2144 5901 2208
rect 5965 2144 5981 2208
rect 6045 2144 6061 2208
rect 6125 2144 6131 2208
rect 5815 2143 6131 2144
rect 8621 2208 8937 2209
rect 8621 2144 8627 2208
rect 8691 2144 8707 2208
rect 8771 2144 8787 2208
rect 8851 2144 8867 2208
rect 8931 2144 8937 2208
rect 8621 2143 8937 2144
rect 11427 2208 11743 2209
rect 11427 2144 11433 2208
rect 11497 2144 11513 2208
rect 11577 2144 11593 2208
rect 11657 2144 11673 2208
rect 11737 2144 11743 2208
rect 11427 2143 11743 2144
<< via3 >>
rect 3015 13084 3079 13088
rect 3015 13028 3019 13084
rect 3019 13028 3075 13084
rect 3075 13028 3079 13084
rect 3015 13024 3079 13028
rect 3095 13084 3159 13088
rect 3095 13028 3099 13084
rect 3099 13028 3155 13084
rect 3155 13028 3159 13084
rect 3095 13024 3159 13028
rect 3175 13084 3239 13088
rect 3175 13028 3179 13084
rect 3179 13028 3235 13084
rect 3235 13028 3239 13084
rect 3175 13024 3239 13028
rect 3255 13084 3319 13088
rect 3255 13028 3259 13084
rect 3259 13028 3315 13084
rect 3315 13028 3319 13084
rect 3255 13024 3319 13028
rect 5821 13084 5885 13088
rect 5821 13028 5825 13084
rect 5825 13028 5881 13084
rect 5881 13028 5885 13084
rect 5821 13024 5885 13028
rect 5901 13084 5965 13088
rect 5901 13028 5905 13084
rect 5905 13028 5961 13084
rect 5961 13028 5965 13084
rect 5901 13024 5965 13028
rect 5981 13084 6045 13088
rect 5981 13028 5985 13084
rect 5985 13028 6041 13084
rect 6041 13028 6045 13084
rect 5981 13024 6045 13028
rect 6061 13084 6125 13088
rect 6061 13028 6065 13084
rect 6065 13028 6121 13084
rect 6121 13028 6125 13084
rect 6061 13024 6125 13028
rect 8627 13084 8691 13088
rect 8627 13028 8631 13084
rect 8631 13028 8687 13084
rect 8687 13028 8691 13084
rect 8627 13024 8691 13028
rect 8707 13084 8771 13088
rect 8707 13028 8711 13084
rect 8711 13028 8767 13084
rect 8767 13028 8771 13084
rect 8707 13024 8771 13028
rect 8787 13084 8851 13088
rect 8787 13028 8791 13084
rect 8791 13028 8847 13084
rect 8847 13028 8851 13084
rect 8787 13024 8851 13028
rect 8867 13084 8931 13088
rect 8867 13028 8871 13084
rect 8871 13028 8927 13084
rect 8927 13028 8931 13084
rect 8867 13024 8931 13028
rect 11433 13084 11497 13088
rect 11433 13028 11437 13084
rect 11437 13028 11493 13084
rect 11493 13028 11497 13084
rect 11433 13024 11497 13028
rect 11513 13084 11577 13088
rect 11513 13028 11517 13084
rect 11517 13028 11573 13084
rect 11573 13028 11577 13084
rect 11513 13024 11577 13028
rect 11593 13084 11657 13088
rect 11593 13028 11597 13084
rect 11597 13028 11653 13084
rect 11653 13028 11657 13084
rect 11593 13024 11657 13028
rect 11673 13084 11737 13088
rect 11673 13028 11677 13084
rect 11677 13028 11733 13084
rect 11733 13028 11737 13084
rect 11673 13024 11737 13028
rect 2355 12540 2419 12544
rect 2355 12484 2359 12540
rect 2359 12484 2415 12540
rect 2415 12484 2419 12540
rect 2355 12480 2419 12484
rect 2435 12540 2499 12544
rect 2435 12484 2439 12540
rect 2439 12484 2495 12540
rect 2495 12484 2499 12540
rect 2435 12480 2499 12484
rect 2515 12540 2579 12544
rect 2515 12484 2519 12540
rect 2519 12484 2575 12540
rect 2575 12484 2579 12540
rect 2515 12480 2579 12484
rect 2595 12540 2659 12544
rect 2595 12484 2599 12540
rect 2599 12484 2655 12540
rect 2655 12484 2659 12540
rect 2595 12480 2659 12484
rect 5161 12540 5225 12544
rect 5161 12484 5165 12540
rect 5165 12484 5221 12540
rect 5221 12484 5225 12540
rect 5161 12480 5225 12484
rect 5241 12540 5305 12544
rect 5241 12484 5245 12540
rect 5245 12484 5301 12540
rect 5301 12484 5305 12540
rect 5241 12480 5305 12484
rect 5321 12540 5385 12544
rect 5321 12484 5325 12540
rect 5325 12484 5381 12540
rect 5381 12484 5385 12540
rect 5321 12480 5385 12484
rect 5401 12540 5465 12544
rect 5401 12484 5405 12540
rect 5405 12484 5461 12540
rect 5461 12484 5465 12540
rect 5401 12480 5465 12484
rect 7967 12540 8031 12544
rect 7967 12484 7971 12540
rect 7971 12484 8027 12540
rect 8027 12484 8031 12540
rect 7967 12480 8031 12484
rect 8047 12540 8111 12544
rect 8047 12484 8051 12540
rect 8051 12484 8107 12540
rect 8107 12484 8111 12540
rect 8047 12480 8111 12484
rect 8127 12540 8191 12544
rect 8127 12484 8131 12540
rect 8131 12484 8187 12540
rect 8187 12484 8191 12540
rect 8127 12480 8191 12484
rect 8207 12540 8271 12544
rect 8207 12484 8211 12540
rect 8211 12484 8267 12540
rect 8267 12484 8271 12540
rect 8207 12480 8271 12484
rect 10773 12540 10837 12544
rect 10773 12484 10777 12540
rect 10777 12484 10833 12540
rect 10833 12484 10837 12540
rect 10773 12480 10837 12484
rect 10853 12540 10917 12544
rect 10853 12484 10857 12540
rect 10857 12484 10913 12540
rect 10913 12484 10917 12540
rect 10853 12480 10917 12484
rect 10933 12540 10997 12544
rect 10933 12484 10937 12540
rect 10937 12484 10993 12540
rect 10993 12484 10997 12540
rect 10933 12480 10997 12484
rect 11013 12540 11077 12544
rect 11013 12484 11017 12540
rect 11017 12484 11073 12540
rect 11073 12484 11077 12540
rect 11013 12480 11077 12484
rect 3015 11996 3079 12000
rect 3015 11940 3019 11996
rect 3019 11940 3075 11996
rect 3075 11940 3079 11996
rect 3015 11936 3079 11940
rect 3095 11996 3159 12000
rect 3095 11940 3099 11996
rect 3099 11940 3155 11996
rect 3155 11940 3159 11996
rect 3095 11936 3159 11940
rect 3175 11996 3239 12000
rect 3175 11940 3179 11996
rect 3179 11940 3235 11996
rect 3235 11940 3239 11996
rect 3175 11936 3239 11940
rect 3255 11996 3319 12000
rect 3255 11940 3259 11996
rect 3259 11940 3315 11996
rect 3315 11940 3319 11996
rect 3255 11936 3319 11940
rect 5821 11996 5885 12000
rect 5821 11940 5825 11996
rect 5825 11940 5881 11996
rect 5881 11940 5885 11996
rect 5821 11936 5885 11940
rect 5901 11996 5965 12000
rect 5901 11940 5905 11996
rect 5905 11940 5961 11996
rect 5961 11940 5965 11996
rect 5901 11936 5965 11940
rect 5981 11996 6045 12000
rect 5981 11940 5985 11996
rect 5985 11940 6041 11996
rect 6041 11940 6045 11996
rect 5981 11936 6045 11940
rect 6061 11996 6125 12000
rect 6061 11940 6065 11996
rect 6065 11940 6121 11996
rect 6121 11940 6125 11996
rect 6061 11936 6125 11940
rect 8627 11996 8691 12000
rect 8627 11940 8631 11996
rect 8631 11940 8687 11996
rect 8687 11940 8691 11996
rect 8627 11936 8691 11940
rect 8707 11996 8771 12000
rect 8707 11940 8711 11996
rect 8711 11940 8767 11996
rect 8767 11940 8771 11996
rect 8707 11936 8771 11940
rect 8787 11996 8851 12000
rect 8787 11940 8791 11996
rect 8791 11940 8847 11996
rect 8847 11940 8851 11996
rect 8787 11936 8851 11940
rect 8867 11996 8931 12000
rect 8867 11940 8871 11996
rect 8871 11940 8927 11996
rect 8927 11940 8931 11996
rect 8867 11936 8931 11940
rect 11433 11996 11497 12000
rect 11433 11940 11437 11996
rect 11437 11940 11493 11996
rect 11493 11940 11497 11996
rect 11433 11936 11497 11940
rect 11513 11996 11577 12000
rect 11513 11940 11517 11996
rect 11517 11940 11573 11996
rect 11573 11940 11577 11996
rect 11513 11936 11577 11940
rect 11593 11996 11657 12000
rect 11593 11940 11597 11996
rect 11597 11940 11653 11996
rect 11653 11940 11657 11996
rect 11593 11936 11657 11940
rect 11673 11996 11737 12000
rect 11673 11940 11677 11996
rect 11677 11940 11733 11996
rect 11733 11940 11737 11996
rect 11673 11936 11737 11940
rect 4108 11596 4172 11660
rect 2355 11452 2419 11456
rect 2355 11396 2359 11452
rect 2359 11396 2415 11452
rect 2415 11396 2419 11452
rect 2355 11392 2419 11396
rect 2435 11452 2499 11456
rect 2435 11396 2439 11452
rect 2439 11396 2495 11452
rect 2495 11396 2499 11452
rect 2435 11392 2499 11396
rect 2515 11452 2579 11456
rect 2515 11396 2519 11452
rect 2519 11396 2575 11452
rect 2575 11396 2579 11452
rect 2515 11392 2579 11396
rect 2595 11452 2659 11456
rect 2595 11396 2599 11452
rect 2599 11396 2655 11452
rect 2655 11396 2659 11452
rect 2595 11392 2659 11396
rect 5161 11452 5225 11456
rect 5161 11396 5165 11452
rect 5165 11396 5221 11452
rect 5221 11396 5225 11452
rect 5161 11392 5225 11396
rect 5241 11452 5305 11456
rect 5241 11396 5245 11452
rect 5245 11396 5301 11452
rect 5301 11396 5305 11452
rect 5241 11392 5305 11396
rect 5321 11452 5385 11456
rect 5321 11396 5325 11452
rect 5325 11396 5381 11452
rect 5381 11396 5385 11452
rect 5321 11392 5385 11396
rect 5401 11452 5465 11456
rect 5401 11396 5405 11452
rect 5405 11396 5461 11452
rect 5461 11396 5465 11452
rect 5401 11392 5465 11396
rect 7967 11452 8031 11456
rect 7967 11396 7971 11452
rect 7971 11396 8027 11452
rect 8027 11396 8031 11452
rect 7967 11392 8031 11396
rect 8047 11452 8111 11456
rect 8047 11396 8051 11452
rect 8051 11396 8107 11452
rect 8107 11396 8111 11452
rect 8047 11392 8111 11396
rect 8127 11452 8191 11456
rect 8127 11396 8131 11452
rect 8131 11396 8187 11452
rect 8187 11396 8191 11452
rect 8127 11392 8191 11396
rect 8207 11452 8271 11456
rect 8207 11396 8211 11452
rect 8211 11396 8267 11452
rect 8267 11396 8271 11452
rect 8207 11392 8271 11396
rect 10773 11452 10837 11456
rect 10773 11396 10777 11452
rect 10777 11396 10833 11452
rect 10833 11396 10837 11452
rect 10773 11392 10837 11396
rect 10853 11452 10917 11456
rect 10853 11396 10857 11452
rect 10857 11396 10913 11452
rect 10913 11396 10917 11452
rect 10853 11392 10917 11396
rect 10933 11452 10997 11456
rect 10933 11396 10937 11452
rect 10937 11396 10993 11452
rect 10993 11396 10997 11452
rect 10933 11392 10997 11396
rect 11013 11452 11077 11456
rect 11013 11396 11017 11452
rect 11017 11396 11073 11452
rect 11073 11396 11077 11452
rect 11013 11392 11077 11396
rect 3015 10908 3079 10912
rect 3015 10852 3019 10908
rect 3019 10852 3075 10908
rect 3075 10852 3079 10908
rect 3015 10848 3079 10852
rect 3095 10908 3159 10912
rect 3095 10852 3099 10908
rect 3099 10852 3155 10908
rect 3155 10852 3159 10908
rect 3095 10848 3159 10852
rect 3175 10908 3239 10912
rect 3175 10852 3179 10908
rect 3179 10852 3235 10908
rect 3235 10852 3239 10908
rect 3175 10848 3239 10852
rect 3255 10908 3319 10912
rect 3255 10852 3259 10908
rect 3259 10852 3315 10908
rect 3315 10852 3319 10908
rect 3255 10848 3319 10852
rect 5821 10908 5885 10912
rect 5821 10852 5825 10908
rect 5825 10852 5881 10908
rect 5881 10852 5885 10908
rect 5821 10848 5885 10852
rect 5901 10908 5965 10912
rect 5901 10852 5905 10908
rect 5905 10852 5961 10908
rect 5961 10852 5965 10908
rect 5901 10848 5965 10852
rect 5981 10908 6045 10912
rect 5981 10852 5985 10908
rect 5985 10852 6041 10908
rect 6041 10852 6045 10908
rect 5981 10848 6045 10852
rect 6061 10908 6125 10912
rect 6061 10852 6065 10908
rect 6065 10852 6121 10908
rect 6121 10852 6125 10908
rect 6061 10848 6125 10852
rect 8627 10908 8691 10912
rect 8627 10852 8631 10908
rect 8631 10852 8687 10908
rect 8687 10852 8691 10908
rect 8627 10848 8691 10852
rect 8707 10908 8771 10912
rect 8707 10852 8711 10908
rect 8711 10852 8767 10908
rect 8767 10852 8771 10908
rect 8707 10848 8771 10852
rect 8787 10908 8851 10912
rect 8787 10852 8791 10908
rect 8791 10852 8847 10908
rect 8847 10852 8851 10908
rect 8787 10848 8851 10852
rect 8867 10908 8931 10912
rect 8867 10852 8871 10908
rect 8871 10852 8927 10908
rect 8927 10852 8931 10908
rect 8867 10848 8931 10852
rect 11433 10908 11497 10912
rect 11433 10852 11437 10908
rect 11437 10852 11493 10908
rect 11493 10852 11497 10908
rect 11433 10848 11497 10852
rect 11513 10908 11577 10912
rect 11513 10852 11517 10908
rect 11517 10852 11573 10908
rect 11573 10852 11577 10908
rect 11513 10848 11577 10852
rect 11593 10908 11657 10912
rect 11593 10852 11597 10908
rect 11597 10852 11653 10908
rect 11653 10852 11657 10908
rect 11593 10848 11657 10852
rect 11673 10908 11737 10912
rect 11673 10852 11677 10908
rect 11677 10852 11733 10908
rect 11733 10852 11737 10908
rect 11673 10848 11737 10852
rect 2355 10364 2419 10368
rect 2355 10308 2359 10364
rect 2359 10308 2415 10364
rect 2415 10308 2419 10364
rect 2355 10304 2419 10308
rect 2435 10364 2499 10368
rect 2435 10308 2439 10364
rect 2439 10308 2495 10364
rect 2495 10308 2499 10364
rect 2435 10304 2499 10308
rect 2515 10364 2579 10368
rect 2515 10308 2519 10364
rect 2519 10308 2575 10364
rect 2575 10308 2579 10364
rect 2515 10304 2579 10308
rect 2595 10364 2659 10368
rect 2595 10308 2599 10364
rect 2599 10308 2655 10364
rect 2655 10308 2659 10364
rect 2595 10304 2659 10308
rect 5161 10364 5225 10368
rect 5161 10308 5165 10364
rect 5165 10308 5221 10364
rect 5221 10308 5225 10364
rect 5161 10304 5225 10308
rect 5241 10364 5305 10368
rect 5241 10308 5245 10364
rect 5245 10308 5301 10364
rect 5301 10308 5305 10364
rect 5241 10304 5305 10308
rect 5321 10364 5385 10368
rect 5321 10308 5325 10364
rect 5325 10308 5381 10364
rect 5381 10308 5385 10364
rect 5321 10304 5385 10308
rect 5401 10364 5465 10368
rect 5401 10308 5405 10364
rect 5405 10308 5461 10364
rect 5461 10308 5465 10364
rect 5401 10304 5465 10308
rect 7967 10364 8031 10368
rect 7967 10308 7971 10364
rect 7971 10308 8027 10364
rect 8027 10308 8031 10364
rect 7967 10304 8031 10308
rect 8047 10364 8111 10368
rect 8047 10308 8051 10364
rect 8051 10308 8107 10364
rect 8107 10308 8111 10364
rect 8047 10304 8111 10308
rect 8127 10364 8191 10368
rect 8127 10308 8131 10364
rect 8131 10308 8187 10364
rect 8187 10308 8191 10364
rect 8127 10304 8191 10308
rect 8207 10364 8271 10368
rect 8207 10308 8211 10364
rect 8211 10308 8267 10364
rect 8267 10308 8271 10364
rect 8207 10304 8271 10308
rect 10773 10364 10837 10368
rect 10773 10308 10777 10364
rect 10777 10308 10833 10364
rect 10833 10308 10837 10364
rect 10773 10304 10837 10308
rect 10853 10364 10917 10368
rect 10853 10308 10857 10364
rect 10857 10308 10913 10364
rect 10913 10308 10917 10364
rect 10853 10304 10917 10308
rect 10933 10364 10997 10368
rect 10933 10308 10937 10364
rect 10937 10308 10993 10364
rect 10993 10308 10997 10364
rect 10933 10304 10997 10308
rect 11013 10364 11077 10368
rect 11013 10308 11017 10364
rect 11017 10308 11073 10364
rect 11073 10308 11077 10364
rect 11013 10304 11077 10308
rect 3015 9820 3079 9824
rect 3015 9764 3019 9820
rect 3019 9764 3075 9820
rect 3075 9764 3079 9820
rect 3015 9760 3079 9764
rect 3095 9820 3159 9824
rect 3095 9764 3099 9820
rect 3099 9764 3155 9820
rect 3155 9764 3159 9820
rect 3095 9760 3159 9764
rect 3175 9820 3239 9824
rect 3175 9764 3179 9820
rect 3179 9764 3235 9820
rect 3235 9764 3239 9820
rect 3175 9760 3239 9764
rect 3255 9820 3319 9824
rect 3255 9764 3259 9820
rect 3259 9764 3315 9820
rect 3315 9764 3319 9820
rect 3255 9760 3319 9764
rect 5821 9820 5885 9824
rect 5821 9764 5825 9820
rect 5825 9764 5881 9820
rect 5881 9764 5885 9820
rect 5821 9760 5885 9764
rect 5901 9820 5965 9824
rect 5901 9764 5905 9820
rect 5905 9764 5961 9820
rect 5961 9764 5965 9820
rect 5901 9760 5965 9764
rect 5981 9820 6045 9824
rect 5981 9764 5985 9820
rect 5985 9764 6041 9820
rect 6041 9764 6045 9820
rect 5981 9760 6045 9764
rect 6061 9820 6125 9824
rect 6061 9764 6065 9820
rect 6065 9764 6121 9820
rect 6121 9764 6125 9820
rect 6061 9760 6125 9764
rect 8627 9820 8691 9824
rect 8627 9764 8631 9820
rect 8631 9764 8687 9820
rect 8687 9764 8691 9820
rect 8627 9760 8691 9764
rect 8707 9820 8771 9824
rect 8707 9764 8711 9820
rect 8711 9764 8767 9820
rect 8767 9764 8771 9820
rect 8707 9760 8771 9764
rect 8787 9820 8851 9824
rect 8787 9764 8791 9820
rect 8791 9764 8847 9820
rect 8847 9764 8851 9820
rect 8787 9760 8851 9764
rect 8867 9820 8931 9824
rect 8867 9764 8871 9820
rect 8871 9764 8927 9820
rect 8927 9764 8931 9820
rect 8867 9760 8931 9764
rect 11433 9820 11497 9824
rect 11433 9764 11437 9820
rect 11437 9764 11493 9820
rect 11493 9764 11497 9820
rect 11433 9760 11497 9764
rect 11513 9820 11577 9824
rect 11513 9764 11517 9820
rect 11517 9764 11573 9820
rect 11573 9764 11577 9820
rect 11513 9760 11577 9764
rect 11593 9820 11657 9824
rect 11593 9764 11597 9820
rect 11597 9764 11653 9820
rect 11653 9764 11657 9820
rect 11593 9760 11657 9764
rect 11673 9820 11737 9824
rect 11673 9764 11677 9820
rect 11677 9764 11733 9820
rect 11733 9764 11737 9820
rect 11673 9760 11737 9764
rect 2355 9276 2419 9280
rect 2355 9220 2359 9276
rect 2359 9220 2415 9276
rect 2415 9220 2419 9276
rect 2355 9216 2419 9220
rect 2435 9276 2499 9280
rect 2435 9220 2439 9276
rect 2439 9220 2495 9276
rect 2495 9220 2499 9276
rect 2435 9216 2499 9220
rect 2515 9276 2579 9280
rect 2515 9220 2519 9276
rect 2519 9220 2575 9276
rect 2575 9220 2579 9276
rect 2515 9216 2579 9220
rect 2595 9276 2659 9280
rect 2595 9220 2599 9276
rect 2599 9220 2655 9276
rect 2655 9220 2659 9276
rect 2595 9216 2659 9220
rect 5161 9276 5225 9280
rect 5161 9220 5165 9276
rect 5165 9220 5221 9276
rect 5221 9220 5225 9276
rect 5161 9216 5225 9220
rect 5241 9276 5305 9280
rect 5241 9220 5245 9276
rect 5245 9220 5301 9276
rect 5301 9220 5305 9276
rect 5241 9216 5305 9220
rect 5321 9276 5385 9280
rect 5321 9220 5325 9276
rect 5325 9220 5381 9276
rect 5381 9220 5385 9276
rect 5321 9216 5385 9220
rect 5401 9276 5465 9280
rect 5401 9220 5405 9276
rect 5405 9220 5461 9276
rect 5461 9220 5465 9276
rect 5401 9216 5465 9220
rect 7967 9276 8031 9280
rect 7967 9220 7971 9276
rect 7971 9220 8027 9276
rect 8027 9220 8031 9276
rect 7967 9216 8031 9220
rect 8047 9276 8111 9280
rect 8047 9220 8051 9276
rect 8051 9220 8107 9276
rect 8107 9220 8111 9276
rect 8047 9216 8111 9220
rect 8127 9276 8191 9280
rect 8127 9220 8131 9276
rect 8131 9220 8187 9276
rect 8187 9220 8191 9276
rect 8127 9216 8191 9220
rect 8207 9276 8271 9280
rect 8207 9220 8211 9276
rect 8211 9220 8267 9276
rect 8267 9220 8271 9276
rect 8207 9216 8271 9220
rect 10773 9276 10837 9280
rect 10773 9220 10777 9276
rect 10777 9220 10833 9276
rect 10833 9220 10837 9276
rect 10773 9216 10837 9220
rect 10853 9276 10917 9280
rect 10853 9220 10857 9276
rect 10857 9220 10913 9276
rect 10913 9220 10917 9276
rect 10853 9216 10917 9220
rect 10933 9276 10997 9280
rect 10933 9220 10937 9276
rect 10937 9220 10993 9276
rect 10993 9220 10997 9276
rect 10933 9216 10997 9220
rect 11013 9276 11077 9280
rect 11013 9220 11017 9276
rect 11017 9220 11073 9276
rect 11073 9220 11077 9276
rect 11013 9216 11077 9220
rect 3015 8732 3079 8736
rect 3015 8676 3019 8732
rect 3019 8676 3075 8732
rect 3075 8676 3079 8732
rect 3015 8672 3079 8676
rect 3095 8732 3159 8736
rect 3095 8676 3099 8732
rect 3099 8676 3155 8732
rect 3155 8676 3159 8732
rect 3095 8672 3159 8676
rect 3175 8732 3239 8736
rect 3175 8676 3179 8732
rect 3179 8676 3235 8732
rect 3235 8676 3239 8732
rect 3175 8672 3239 8676
rect 3255 8732 3319 8736
rect 3255 8676 3259 8732
rect 3259 8676 3315 8732
rect 3315 8676 3319 8732
rect 3255 8672 3319 8676
rect 5821 8732 5885 8736
rect 5821 8676 5825 8732
rect 5825 8676 5881 8732
rect 5881 8676 5885 8732
rect 5821 8672 5885 8676
rect 5901 8732 5965 8736
rect 5901 8676 5905 8732
rect 5905 8676 5961 8732
rect 5961 8676 5965 8732
rect 5901 8672 5965 8676
rect 5981 8732 6045 8736
rect 5981 8676 5985 8732
rect 5985 8676 6041 8732
rect 6041 8676 6045 8732
rect 5981 8672 6045 8676
rect 6061 8732 6125 8736
rect 6061 8676 6065 8732
rect 6065 8676 6121 8732
rect 6121 8676 6125 8732
rect 6061 8672 6125 8676
rect 8627 8732 8691 8736
rect 8627 8676 8631 8732
rect 8631 8676 8687 8732
rect 8687 8676 8691 8732
rect 8627 8672 8691 8676
rect 8707 8732 8771 8736
rect 8707 8676 8711 8732
rect 8711 8676 8767 8732
rect 8767 8676 8771 8732
rect 8707 8672 8771 8676
rect 8787 8732 8851 8736
rect 8787 8676 8791 8732
rect 8791 8676 8847 8732
rect 8847 8676 8851 8732
rect 8787 8672 8851 8676
rect 8867 8732 8931 8736
rect 8867 8676 8871 8732
rect 8871 8676 8927 8732
rect 8927 8676 8931 8732
rect 8867 8672 8931 8676
rect 11433 8732 11497 8736
rect 11433 8676 11437 8732
rect 11437 8676 11493 8732
rect 11493 8676 11497 8732
rect 11433 8672 11497 8676
rect 11513 8732 11577 8736
rect 11513 8676 11517 8732
rect 11517 8676 11573 8732
rect 11573 8676 11577 8732
rect 11513 8672 11577 8676
rect 11593 8732 11657 8736
rect 11593 8676 11597 8732
rect 11597 8676 11653 8732
rect 11653 8676 11657 8732
rect 11593 8672 11657 8676
rect 11673 8732 11737 8736
rect 11673 8676 11677 8732
rect 11677 8676 11733 8732
rect 11733 8676 11737 8732
rect 11673 8672 11737 8676
rect 4108 8196 4172 8260
rect 2355 8188 2419 8192
rect 2355 8132 2359 8188
rect 2359 8132 2415 8188
rect 2415 8132 2419 8188
rect 2355 8128 2419 8132
rect 2435 8188 2499 8192
rect 2435 8132 2439 8188
rect 2439 8132 2495 8188
rect 2495 8132 2499 8188
rect 2435 8128 2499 8132
rect 2515 8188 2579 8192
rect 2515 8132 2519 8188
rect 2519 8132 2575 8188
rect 2575 8132 2579 8188
rect 2515 8128 2579 8132
rect 2595 8188 2659 8192
rect 2595 8132 2599 8188
rect 2599 8132 2655 8188
rect 2655 8132 2659 8188
rect 2595 8128 2659 8132
rect 5161 8188 5225 8192
rect 5161 8132 5165 8188
rect 5165 8132 5221 8188
rect 5221 8132 5225 8188
rect 5161 8128 5225 8132
rect 5241 8188 5305 8192
rect 5241 8132 5245 8188
rect 5245 8132 5301 8188
rect 5301 8132 5305 8188
rect 5241 8128 5305 8132
rect 5321 8188 5385 8192
rect 5321 8132 5325 8188
rect 5325 8132 5381 8188
rect 5381 8132 5385 8188
rect 5321 8128 5385 8132
rect 5401 8188 5465 8192
rect 5401 8132 5405 8188
rect 5405 8132 5461 8188
rect 5461 8132 5465 8188
rect 5401 8128 5465 8132
rect 7967 8188 8031 8192
rect 7967 8132 7971 8188
rect 7971 8132 8027 8188
rect 8027 8132 8031 8188
rect 7967 8128 8031 8132
rect 8047 8188 8111 8192
rect 8047 8132 8051 8188
rect 8051 8132 8107 8188
rect 8107 8132 8111 8188
rect 8047 8128 8111 8132
rect 8127 8188 8191 8192
rect 8127 8132 8131 8188
rect 8131 8132 8187 8188
rect 8187 8132 8191 8188
rect 8127 8128 8191 8132
rect 8207 8188 8271 8192
rect 8207 8132 8211 8188
rect 8211 8132 8267 8188
rect 8267 8132 8271 8188
rect 8207 8128 8271 8132
rect 10773 8188 10837 8192
rect 10773 8132 10777 8188
rect 10777 8132 10833 8188
rect 10833 8132 10837 8188
rect 10773 8128 10837 8132
rect 10853 8188 10917 8192
rect 10853 8132 10857 8188
rect 10857 8132 10913 8188
rect 10913 8132 10917 8188
rect 10853 8128 10917 8132
rect 10933 8188 10997 8192
rect 10933 8132 10937 8188
rect 10937 8132 10993 8188
rect 10993 8132 10997 8188
rect 10933 8128 10997 8132
rect 11013 8188 11077 8192
rect 11013 8132 11017 8188
rect 11017 8132 11073 8188
rect 11073 8132 11077 8188
rect 11013 8128 11077 8132
rect 3015 7644 3079 7648
rect 3015 7588 3019 7644
rect 3019 7588 3075 7644
rect 3075 7588 3079 7644
rect 3015 7584 3079 7588
rect 3095 7644 3159 7648
rect 3095 7588 3099 7644
rect 3099 7588 3155 7644
rect 3155 7588 3159 7644
rect 3095 7584 3159 7588
rect 3175 7644 3239 7648
rect 3175 7588 3179 7644
rect 3179 7588 3235 7644
rect 3235 7588 3239 7644
rect 3175 7584 3239 7588
rect 3255 7644 3319 7648
rect 3255 7588 3259 7644
rect 3259 7588 3315 7644
rect 3315 7588 3319 7644
rect 3255 7584 3319 7588
rect 5821 7644 5885 7648
rect 5821 7588 5825 7644
rect 5825 7588 5881 7644
rect 5881 7588 5885 7644
rect 5821 7584 5885 7588
rect 5901 7644 5965 7648
rect 5901 7588 5905 7644
rect 5905 7588 5961 7644
rect 5961 7588 5965 7644
rect 5901 7584 5965 7588
rect 5981 7644 6045 7648
rect 5981 7588 5985 7644
rect 5985 7588 6041 7644
rect 6041 7588 6045 7644
rect 5981 7584 6045 7588
rect 6061 7644 6125 7648
rect 6061 7588 6065 7644
rect 6065 7588 6121 7644
rect 6121 7588 6125 7644
rect 6061 7584 6125 7588
rect 8627 7644 8691 7648
rect 8627 7588 8631 7644
rect 8631 7588 8687 7644
rect 8687 7588 8691 7644
rect 8627 7584 8691 7588
rect 8707 7644 8771 7648
rect 8707 7588 8711 7644
rect 8711 7588 8767 7644
rect 8767 7588 8771 7644
rect 8707 7584 8771 7588
rect 8787 7644 8851 7648
rect 8787 7588 8791 7644
rect 8791 7588 8847 7644
rect 8847 7588 8851 7644
rect 8787 7584 8851 7588
rect 8867 7644 8931 7648
rect 8867 7588 8871 7644
rect 8871 7588 8927 7644
rect 8927 7588 8931 7644
rect 8867 7584 8931 7588
rect 11433 7644 11497 7648
rect 11433 7588 11437 7644
rect 11437 7588 11493 7644
rect 11493 7588 11497 7644
rect 11433 7584 11497 7588
rect 11513 7644 11577 7648
rect 11513 7588 11517 7644
rect 11517 7588 11573 7644
rect 11573 7588 11577 7644
rect 11513 7584 11577 7588
rect 11593 7644 11657 7648
rect 11593 7588 11597 7644
rect 11597 7588 11653 7644
rect 11653 7588 11657 7644
rect 11593 7584 11657 7588
rect 11673 7644 11737 7648
rect 11673 7588 11677 7644
rect 11677 7588 11733 7644
rect 11733 7588 11737 7644
rect 11673 7584 11737 7588
rect 2355 7100 2419 7104
rect 2355 7044 2359 7100
rect 2359 7044 2415 7100
rect 2415 7044 2419 7100
rect 2355 7040 2419 7044
rect 2435 7100 2499 7104
rect 2435 7044 2439 7100
rect 2439 7044 2495 7100
rect 2495 7044 2499 7100
rect 2435 7040 2499 7044
rect 2515 7100 2579 7104
rect 2515 7044 2519 7100
rect 2519 7044 2575 7100
rect 2575 7044 2579 7100
rect 2515 7040 2579 7044
rect 2595 7100 2659 7104
rect 2595 7044 2599 7100
rect 2599 7044 2655 7100
rect 2655 7044 2659 7100
rect 2595 7040 2659 7044
rect 5161 7100 5225 7104
rect 5161 7044 5165 7100
rect 5165 7044 5221 7100
rect 5221 7044 5225 7100
rect 5161 7040 5225 7044
rect 5241 7100 5305 7104
rect 5241 7044 5245 7100
rect 5245 7044 5301 7100
rect 5301 7044 5305 7100
rect 5241 7040 5305 7044
rect 5321 7100 5385 7104
rect 5321 7044 5325 7100
rect 5325 7044 5381 7100
rect 5381 7044 5385 7100
rect 5321 7040 5385 7044
rect 5401 7100 5465 7104
rect 5401 7044 5405 7100
rect 5405 7044 5461 7100
rect 5461 7044 5465 7100
rect 5401 7040 5465 7044
rect 7967 7100 8031 7104
rect 7967 7044 7971 7100
rect 7971 7044 8027 7100
rect 8027 7044 8031 7100
rect 7967 7040 8031 7044
rect 8047 7100 8111 7104
rect 8047 7044 8051 7100
rect 8051 7044 8107 7100
rect 8107 7044 8111 7100
rect 8047 7040 8111 7044
rect 8127 7100 8191 7104
rect 8127 7044 8131 7100
rect 8131 7044 8187 7100
rect 8187 7044 8191 7100
rect 8127 7040 8191 7044
rect 8207 7100 8271 7104
rect 8207 7044 8211 7100
rect 8211 7044 8267 7100
rect 8267 7044 8271 7100
rect 8207 7040 8271 7044
rect 10773 7100 10837 7104
rect 10773 7044 10777 7100
rect 10777 7044 10833 7100
rect 10833 7044 10837 7100
rect 10773 7040 10837 7044
rect 10853 7100 10917 7104
rect 10853 7044 10857 7100
rect 10857 7044 10913 7100
rect 10913 7044 10917 7100
rect 10853 7040 10917 7044
rect 10933 7100 10997 7104
rect 10933 7044 10937 7100
rect 10937 7044 10993 7100
rect 10993 7044 10997 7100
rect 10933 7040 10997 7044
rect 11013 7100 11077 7104
rect 11013 7044 11017 7100
rect 11017 7044 11073 7100
rect 11073 7044 11077 7100
rect 11013 7040 11077 7044
rect 3015 6556 3079 6560
rect 3015 6500 3019 6556
rect 3019 6500 3075 6556
rect 3075 6500 3079 6556
rect 3015 6496 3079 6500
rect 3095 6556 3159 6560
rect 3095 6500 3099 6556
rect 3099 6500 3155 6556
rect 3155 6500 3159 6556
rect 3095 6496 3159 6500
rect 3175 6556 3239 6560
rect 3175 6500 3179 6556
rect 3179 6500 3235 6556
rect 3235 6500 3239 6556
rect 3175 6496 3239 6500
rect 3255 6556 3319 6560
rect 3255 6500 3259 6556
rect 3259 6500 3315 6556
rect 3315 6500 3319 6556
rect 3255 6496 3319 6500
rect 5821 6556 5885 6560
rect 5821 6500 5825 6556
rect 5825 6500 5881 6556
rect 5881 6500 5885 6556
rect 5821 6496 5885 6500
rect 5901 6556 5965 6560
rect 5901 6500 5905 6556
rect 5905 6500 5961 6556
rect 5961 6500 5965 6556
rect 5901 6496 5965 6500
rect 5981 6556 6045 6560
rect 5981 6500 5985 6556
rect 5985 6500 6041 6556
rect 6041 6500 6045 6556
rect 5981 6496 6045 6500
rect 6061 6556 6125 6560
rect 6061 6500 6065 6556
rect 6065 6500 6121 6556
rect 6121 6500 6125 6556
rect 6061 6496 6125 6500
rect 8627 6556 8691 6560
rect 8627 6500 8631 6556
rect 8631 6500 8687 6556
rect 8687 6500 8691 6556
rect 8627 6496 8691 6500
rect 8707 6556 8771 6560
rect 8707 6500 8711 6556
rect 8711 6500 8767 6556
rect 8767 6500 8771 6556
rect 8707 6496 8771 6500
rect 8787 6556 8851 6560
rect 8787 6500 8791 6556
rect 8791 6500 8847 6556
rect 8847 6500 8851 6556
rect 8787 6496 8851 6500
rect 8867 6556 8931 6560
rect 8867 6500 8871 6556
rect 8871 6500 8927 6556
rect 8927 6500 8931 6556
rect 8867 6496 8931 6500
rect 11433 6556 11497 6560
rect 11433 6500 11437 6556
rect 11437 6500 11493 6556
rect 11493 6500 11497 6556
rect 11433 6496 11497 6500
rect 11513 6556 11577 6560
rect 11513 6500 11517 6556
rect 11517 6500 11573 6556
rect 11573 6500 11577 6556
rect 11513 6496 11577 6500
rect 11593 6556 11657 6560
rect 11593 6500 11597 6556
rect 11597 6500 11653 6556
rect 11653 6500 11657 6556
rect 11593 6496 11657 6500
rect 11673 6556 11737 6560
rect 11673 6500 11677 6556
rect 11677 6500 11733 6556
rect 11733 6500 11737 6556
rect 11673 6496 11737 6500
rect 2355 6012 2419 6016
rect 2355 5956 2359 6012
rect 2359 5956 2415 6012
rect 2415 5956 2419 6012
rect 2355 5952 2419 5956
rect 2435 6012 2499 6016
rect 2435 5956 2439 6012
rect 2439 5956 2495 6012
rect 2495 5956 2499 6012
rect 2435 5952 2499 5956
rect 2515 6012 2579 6016
rect 2515 5956 2519 6012
rect 2519 5956 2575 6012
rect 2575 5956 2579 6012
rect 2515 5952 2579 5956
rect 2595 6012 2659 6016
rect 2595 5956 2599 6012
rect 2599 5956 2655 6012
rect 2655 5956 2659 6012
rect 2595 5952 2659 5956
rect 5161 6012 5225 6016
rect 5161 5956 5165 6012
rect 5165 5956 5221 6012
rect 5221 5956 5225 6012
rect 5161 5952 5225 5956
rect 5241 6012 5305 6016
rect 5241 5956 5245 6012
rect 5245 5956 5301 6012
rect 5301 5956 5305 6012
rect 5241 5952 5305 5956
rect 5321 6012 5385 6016
rect 5321 5956 5325 6012
rect 5325 5956 5381 6012
rect 5381 5956 5385 6012
rect 5321 5952 5385 5956
rect 5401 6012 5465 6016
rect 5401 5956 5405 6012
rect 5405 5956 5461 6012
rect 5461 5956 5465 6012
rect 5401 5952 5465 5956
rect 7967 6012 8031 6016
rect 7967 5956 7971 6012
rect 7971 5956 8027 6012
rect 8027 5956 8031 6012
rect 7967 5952 8031 5956
rect 8047 6012 8111 6016
rect 8047 5956 8051 6012
rect 8051 5956 8107 6012
rect 8107 5956 8111 6012
rect 8047 5952 8111 5956
rect 8127 6012 8191 6016
rect 8127 5956 8131 6012
rect 8131 5956 8187 6012
rect 8187 5956 8191 6012
rect 8127 5952 8191 5956
rect 8207 6012 8271 6016
rect 8207 5956 8211 6012
rect 8211 5956 8267 6012
rect 8267 5956 8271 6012
rect 8207 5952 8271 5956
rect 10773 6012 10837 6016
rect 10773 5956 10777 6012
rect 10777 5956 10833 6012
rect 10833 5956 10837 6012
rect 10773 5952 10837 5956
rect 10853 6012 10917 6016
rect 10853 5956 10857 6012
rect 10857 5956 10913 6012
rect 10913 5956 10917 6012
rect 10853 5952 10917 5956
rect 10933 6012 10997 6016
rect 10933 5956 10937 6012
rect 10937 5956 10993 6012
rect 10993 5956 10997 6012
rect 10933 5952 10997 5956
rect 11013 6012 11077 6016
rect 11013 5956 11017 6012
rect 11017 5956 11073 6012
rect 11073 5956 11077 6012
rect 11013 5952 11077 5956
rect 3015 5468 3079 5472
rect 3015 5412 3019 5468
rect 3019 5412 3075 5468
rect 3075 5412 3079 5468
rect 3015 5408 3079 5412
rect 3095 5468 3159 5472
rect 3095 5412 3099 5468
rect 3099 5412 3155 5468
rect 3155 5412 3159 5468
rect 3095 5408 3159 5412
rect 3175 5468 3239 5472
rect 3175 5412 3179 5468
rect 3179 5412 3235 5468
rect 3235 5412 3239 5468
rect 3175 5408 3239 5412
rect 3255 5468 3319 5472
rect 3255 5412 3259 5468
rect 3259 5412 3315 5468
rect 3315 5412 3319 5468
rect 3255 5408 3319 5412
rect 5821 5468 5885 5472
rect 5821 5412 5825 5468
rect 5825 5412 5881 5468
rect 5881 5412 5885 5468
rect 5821 5408 5885 5412
rect 5901 5468 5965 5472
rect 5901 5412 5905 5468
rect 5905 5412 5961 5468
rect 5961 5412 5965 5468
rect 5901 5408 5965 5412
rect 5981 5468 6045 5472
rect 5981 5412 5985 5468
rect 5985 5412 6041 5468
rect 6041 5412 6045 5468
rect 5981 5408 6045 5412
rect 6061 5468 6125 5472
rect 6061 5412 6065 5468
rect 6065 5412 6121 5468
rect 6121 5412 6125 5468
rect 6061 5408 6125 5412
rect 8627 5468 8691 5472
rect 8627 5412 8631 5468
rect 8631 5412 8687 5468
rect 8687 5412 8691 5468
rect 8627 5408 8691 5412
rect 8707 5468 8771 5472
rect 8707 5412 8711 5468
rect 8711 5412 8767 5468
rect 8767 5412 8771 5468
rect 8707 5408 8771 5412
rect 8787 5468 8851 5472
rect 8787 5412 8791 5468
rect 8791 5412 8847 5468
rect 8847 5412 8851 5468
rect 8787 5408 8851 5412
rect 8867 5468 8931 5472
rect 8867 5412 8871 5468
rect 8871 5412 8927 5468
rect 8927 5412 8931 5468
rect 8867 5408 8931 5412
rect 11433 5468 11497 5472
rect 11433 5412 11437 5468
rect 11437 5412 11493 5468
rect 11493 5412 11497 5468
rect 11433 5408 11497 5412
rect 11513 5468 11577 5472
rect 11513 5412 11517 5468
rect 11517 5412 11573 5468
rect 11573 5412 11577 5468
rect 11513 5408 11577 5412
rect 11593 5468 11657 5472
rect 11593 5412 11597 5468
rect 11597 5412 11653 5468
rect 11653 5412 11657 5468
rect 11593 5408 11657 5412
rect 11673 5468 11737 5472
rect 11673 5412 11677 5468
rect 11677 5412 11733 5468
rect 11733 5412 11737 5468
rect 11673 5408 11737 5412
rect 2355 4924 2419 4928
rect 2355 4868 2359 4924
rect 2359 4868 2415 4924
rect 2415 4868 2419 4924
rect 2355 4864 2419 4868
rect 2435 4924 2499 4928
rect 2435 4868 2439 4924
rect 2439 4868 2495 4924
rect 2495 4868 2499 4924
rect 2435 4864 2499 4868
rect 2515 4924 2579 4928
rect 2515 4868 2519 4924
rect 2519 4868 2575 4924
rect 2575 4868 2579 4924
rect 2515 4864 2579 4868
rect 2595 4924 2659 4928
rect 2595 4868 2599 4924
rect 2599 4868 2655 4924
rect 2655 4868 2659 4924
rect 2595 4864 2659 4868
rect 5161 4924 5225 4928
rect 5161 4868 5165 4924
rect 5165 4868 5221 4924
rect 5221 4868 5225 4924
rect 5161 4864 5225 4868
rect 5241 4924 5305 4928
rect 5241 4868 5245 4924
rect 5245 4868 5301 4924
rect 5301 4868 5305 4924
rect 5241 4864 5305 4868
rect 5321 4924 5385 4928
rect 5321 4868 5325 4924
rect 5325 4868 5381 4924
rect 5381 4868 5385 4924
rect 5321 4864 5385 4868
rect 5401 4924 5465 4928
rect 5401 4868 5405 4924
rect 5405 4868 5461 4924
rect 5461 4868 5465 4924
rect 5401 4864 5465 4868
rect 7967 4924 8031 4928
rect 7967 4868 7971 4924
rect 7971 4868 8027 4924
rect 8027 4868 8031 4924
rect 7967 4864 8031 4868
rect 8047 4924 8111 4928
rect 8047 4868 8051 4924
rect 8051 4868 8107 4924
rect 8107 4868 8111 4924
rect 8047 4864 8111 4868
rect 8127 4924 8191 4928
rect 8127 4868 8131 4924
rect 8131 4868 8187 4924
rect 8187 4868 8191 4924
rect 8127 4864 8191 4868
rect 8207 4924 8271 4928
rect 8207 4868 8211 4924
rect 8211 4868 8267 4924
rect 8267 4868 8271 4924
rect 8207 4864 8271 4868
rect 10773 4924 10837 4928
rect 10773 4868 10777 4924
rect 10777 4868 10833 4924
rect 10833 4868 10837 4924
rect 10773 4864 10837 4868
rect 10853 4924 10917 4928
rect 10853 4868 10857 4924
rect 10857 4868 10913 4924
rect 10913 4868 10917 4924
rect 10853 4864 10917 4868
rect 10933 4924 10997 4928
rect 10933 4868 10937 4924
rect 10937 4868 10993 4924
rect 10993 4868 10997 4924
rect 10933 4864 10997 4868
rect 11013 4924 11077 4928
rect 11013 4868 11017 4924
rect 11017 4868 11073 4924
rect 11073 4868 11077 4924
rect 11013 4864 11077 4868
rect 3015 4380 3079 4384
rect 3015 4324 3019 4380
rect 3019 4324 3075 4380
rect 3075 4324 3079 4380
rect 3015 4320 3079 4324
rect 3095 4380 3159 4384
rect 3095 4324 3099 4380
rect 3099 4324 3155 4380
rect 3155 4324 3159 4380
rect 3095 4320 3159 4324
rect 3175 4380 3239 4384
rect 3175 4324 3179 4380
rect 3179 4324 3235 4380
rect 3235 4324 3239 4380
rect 3175 4320 3239 4324
rect 3255 4380 3319 4384
rect 3255 4324 3259 4380
rect 3259 4324 3315 4380
rect 3315 4324 3319 4380
rect 3255 4320 3319 4324
rect 5821 4380 5885 4384
rect 5821 4324 5825 4380
rect 5825 4324 5881 4380
rect 5881 4324 5885 4380
rect 5821 4320 5885 4324
rect 5901 4380 5965 4384
rect 5901 4324 5905 4380
rect 5905 4324 5961 4380
rect 5961 4324 5965 4380
rect 5901 4320 5965 4324
rect 5981 4380 6045 4384
rect 5981 4324 5985 4380
rect 5985 4324 6041 4380
rect 6041 4324 6045 4380
rect 5981 4320 6045 4324
rect 6061 4380 6125 4384
rect 6061 4324 6065 4380
rect 6065 4324 6121 4380
rect 6121 4324 6125 4380
rect 6061 4320 6125 4324
rect 8627 4380 8691 4384
rect 8627 4324 8631 4380
rect 8631 4324 8687 4380
rect 8687 4324 8691 4380
rect 8627 4320 8691 4324
rect 8707 4380 8771 4384
rect 8707 4324 8711 4380
rect 8711 4324 8767 4380
rect 8767 4324 8771 4380
rect 8707 4320 8771 4324
rect 8787 4380 8851 4384
rect 8787 4324 8791 4380
rect 8791 4324 8847 4380
rect 8847 4324 8851 4380
rect 8787 4320 8851 4324
rect 8867 4380 8931 4384
rect 8867 4324 8871 4380
rect 8871 4324 8927 4380
rect 8927 4324 8931 4380
rect 8867 4320 8931 4324
rect 11433 4380 11497 4384
rect 11433 4324 11437 4380
rect 11437 4324 11493 4380
rect 11493 4324 11497 4380
rect 11433 4320 11497 4324
rect 11513 4380 11577 4384
rect 11513 4324 11517 4380
rect 11517 4324 11573 4380
rect 11573 4324 11577 4380
rect 11513 4320 11577 4324
rect 11593 4380 11657 4384
rect 11593 4324 11597 4380
rect 11597 4324 11653 4380
rect 11653 4324 11657 4380
rect 11593 4320 11657 4324
rect 11673 4380 11737 4384
rect 11673 4324 11677 4380
rect 11677 4324 11733 4380
rect 11733 4324 11737 4380
rect 11673 4320 11737 4324
rect 2355 3836 2419 3840
rect 2355 3780 2359 3836
rect 2359 3780 2415 3836
rect 2415 3780 2419 3836
rect 2355 3776 2419 3780
rect 2435 3836 2499 3840
rect 2435 3780 2439 3836
rect 2439 3780 2495 3836
rect 2495 3780 2499 3836
rect 2435 3776 2499 3780
rect 2515 3836 2579 3840
rect 2515 3780 2519 3836
rect 2519 3780 2575 3836
rect 2575 3780 2579 3836
rect 2515 3776 2579 3780
rect 2595 3836 2659 3840
rect 2595 3780 2599 3836
rect 2599 3780 2655 3836
rect 2655 3780 2659 3836
rect 2595 3776 2659 3780
rect 5161 3836 5225 3840
rect 5161 3780 5165 3836
rect 5165 3780 5221 3836
rect 5221 3780 5225 3836
rect 5161 3776 5225 3780
rect 5241 3836 5305 3840
rect 5241 3780 5245 3836
rect 5245 3780 5301 3836
rect 5301 3780 5305 3836
rect 5241 3776 5305 3780
rect 5321 3836 5385 3840
rect 5321 3780 5325 3836
rect 5325 3780 5381 3836
rect 5381 3780 5385 3836
rect 5321 3776 5385 3780
rect 5401 3836 5465 3840
rect 5401 3780 5405 3836
rect 5405 3780 5461 3836
rect 5461 3780 5465 3836
rect 5401 3776 5465 3780
rect 7967 3836 8031 3840
rect 7967 3780 7971 3836
rect 7971 3780 8027 3836
rect 8027 3780 8031 3836
rect 7967 3776 8031 3780
rect 8047 3836 8111 3840
rect 8047 3780 8051 3836
rect 8051 3780 8107 3836
rect 8107 3780 8111 3836
rect 8047 3776 8111 3780
rect 8127 3836 8191 3840
rect 8127 3780 8131 3836
rect 8131 3780 8187 3836
rect 8187 3780 8191 3836
rect 8127 3776 8191 3780
rect 8207 3836 8271 3840
rect 8207 3780 8211 3836
rect 8211 3780 8267 3836
rect 8267 3780 8271 3836
rect 8207 3776 8271 3780
rect 10773 3836 10837 3840
rect 10773 3780 10777 3836
rect 10777 3780 10833 3836
rect 10833 3780 10837 3836
rect 10773 3776 10837 3780
rect 10853 3836 10917 3840
rect 10853 3780 10857 3836
rect 10857 3780 10913 3836
rect 10913 3780 10917 3836
rect 10853 3776 10917 3780
rect 10933 3836 10997 3840
rect 10933 3780 10937 3836
rect 10937 3780 10993 3836
rect 10993 3780 10997 3836
rect 10933 3776 10997 3780
rect 11013 3836 11077 3840
rect 11013 3780 11017 3836
rect 11017 3780 11073 3836
rect 11073 3780 11077 3836
rect 11013 3776 11077 3780
rect 3015 3292 3079 3296
rect 3015 3236 3019 3292
rect 3019 3236 3075 3292
rect 3075 3236 3079 3292
rect 3015 3232 3079 3236
rect 3095 3292 3159 3296
rect 3095 3236 3099 3292
rect 3099 3236 3155 3292
rect 3155 3236 3159 3292
rect 3095 3232 3159 3236
rect 3175 3292 3239 3296
rect 3175 3236 3179 3292
rect 3179 3236 3235 3292
rect 3235 3236 3239 3292
rect 3175 3232 3239 3236
rect 3255 3292 3319 3296
rect 3255 3236 3259 3292
rect 3259 3236 3315 3292
rect 3315 3236 3319 3292
rect 3255 3232 3319 3236
rect 5821 3292 5885 3296
rect 5821 3236 5825 3292
rect 5825 3236 5881 3292
rect 5881 3236 5885 3292
rect 5821 3232 5885 3236
rect 5901 3292 5965 3296
rect 5901 3236 5905 3292
rect 5905 3236 5961 3292
rect 5961 3236 5965 3292
rect 5901 3232 5965 3236
rect 5981 3292 6045 3296
rect 5981 3236 5985 3292
rect 5985 3236 6041 3292
rect 6041 3236 6045 3292
rect 5981 3232 6045 3236
rect 6061 3292 6125 3296
rect 6061 3236 6065 3292
rect 6065 3236 6121 3292
rect 6121 3236 6125 3292
rect 6061 3232 6125 3236
rect 8627 3292 8691 3296
rect 8627 3236 8631 3292
rect 8631 3236 8687 3292
rect 8687 3236 8691 3292
rect 8627 3232 8691 3236
rect 8707 3292 8771 3296
rect 8707 3236 8711 3292
rect 8711 3236 8767 3292
rect 8767 3236 8771 3292
rect 8707 3232 8771 3236
rect 8787 3292 8851 3296
rect 8787 3236 8791 3292
rect 8791 3236 8847 3292
rect 8847 3236 8851 3292
rect 8787 3232 8851 3236
rect 8867 3292 8931 3296
rect 8867 3236 8871 3292
rect 8871 3236 8927 3292
rect 8927 3236 8931 3292
rect 8867 3232 8931 3236
rect 11433 3292 11497 3296
rect 11433 3236 11437 3292
rect 11437 3236 11493 3292
rect 11493 3236 11497 3292
rect 11433 3232 11497 3236
rect 11513 3292 11577 3296
rect 11513 3236 11517 3292
rect 11517 3236 11573 3292
rect 11573 3236 11577 3292
rect 11513 3232 11577 3236
rect 11593 3292 11657 3296
rect 11593 3236 11597 3292
rect 11597 3236 11653 3292
rect 11653 3236 11657 3292
rect 11593 3232 11657 3236
rect 11673 3292 11737 3296
rect 11673 3236 11677 3292
rect 11677 3236 11733 3292
rect 11733 3236 11737 3292
rect 11673 3232 11737 3236
rect 2355 2748 2419 2752
rect 2355 2692 2359 2748
rect 2359 2692 2415 2748
rect 2415 2692 2419 2748
rect 2355 2688 2419 2692
rect 2435 2748 2499 2752
rect 2435 2692 2439 2748
rect 2439 2692 2495 2748
rect 2495 2692 2499 2748
rect 2435 2688 2499 2692
rect 2515 2748 2579 2752
rect 2515 2692 2519 2748
rect 2519 2692 2575 2748
rect 2575 2692 2579 2748
rect 2515 2688 2579 2692
rect 2595 2748 2659 2752
rect 2595 2692 2599 2748
rect 2599 2692 2655 2748
rect 2655 2692 2659 2748
rect 2595 2688 2659 2692
rect 5161 2748 5225 2752
rect 5161 2692 5165 2748
rect 5165 2692 5221 2748
rect 5221 2692 5225 2748
rect 5161 2688 5225 2692
rect 5241 2748 5305 2752
rect 5241 2692 5245 2748
rect 5245 2692 5301 2748
rect 5301 2692 5305 2748
rect 5241 2688 5305 2692
rect 5321 2748 5385 2752
rect 5321 2692 5325 2748
rect 5325 2692 5381 2748
rect 5381 2692 5385 2748
rect 5321 2688 5385 2692
rect 5401 2748 5465 2752
rect 5401 2692 5405 2748
rect 5405 2692 5461 2748
rect 5461 2692 5465 2748
rect 5401 2688 5465 2692
rect 7967 2748 8031 2752
rect 7967 2692 7971 2748
rect 7971 2692 8027 2748
rect 8027 2692 8031 2748
rect 7967 2688 8031 2692
rect 8047 2748 8111 2752
rect 8047 2692 8051 2748
rect 8051 2692 8107 2748
rect 8107 2692 8111 2748
rect 8047 2688 8111 2692
rect 8127 2748 8191 2752
rect 8127 2692 8131 2748
rect 8131 2692 8187 2748
rect 8187 2692 8191 2748
rect 8127 2688 8191 2692
rect 8207 2748 8271 2752
rect 8207 2692 8211 2748
rect 8211 2692 8267 2748
rect 8267 2692 8271 2748
rect 8207 2688 8271 2692
rect 10773 2748 10837 2752
rect 10773 2692 10777 2748
rect 10777 2692 10833 2748
rect 10833 2692 10837 2748
rect 10773 2688 10837 2692
rect 10853 2748 10917 2752
rect 10853 2692 10857 2748
rect 10857 2692 10913 2748
rect 10913 2692 10917 2748
rect 10853 2688 10917 2692
rect 10933 2748 10997 2752
rect 10933 2692 10937 2748
rect 10937 2692 10993 2748
rect 10993 2692 10997 2748
rect 10933 2688 10997 2692
rect 11013 2748 11077 2752
rect 11013 2692 11017 2748
rect 11017 2692 11073 2748
rect 11073 2692 11077 2748
rect 11013 2688 11077 2692
rect 3015 2204 3079 2208
rect 3015 2148 3019 2204
rect 3019 2148 3075 2204
rect 3075 2148 3079 2204
rect 3015 2144 3079 2148
rect 3095 2204 3159 2208
rect 3095 2148 3099 2204
rect 3099 2148 3155 2204
rect 3155 2148 3159 2204
rect 3095 2144 3159 2148
rect 3175 2204 3239 2208
rect 3175 2148 3179 2204
rect 3179 2148 3235 2204
rect 3235 2148 3239 2204
rect 3175 2144 3239 2148
rect 3255 2204 3319 2208
rect 3255 2148 3259 2204
rect 3259 2148 3315 2204
rect 3315 2148 3319 2204
rect 3255 2144 3319 2148
rect 5821 2204 5885 2208
rect 5821 2148 5825 2204
rect 5825 2148 5881 2204
rect 5881 2148 5885 2204
rect 5821 2144 5885 2148
rect 5901 2204 5965 2208
rect 5901 2148 5905 2204
rect 5905 2148 5961 2204
rect 5961 2148 5965 2204
rect 5901 2144 5965 2148
rect 5981 2204 6045 2208
rect 5981 2148 5985 2204
rect 5985 2148 6041 2204
rect 6041 2148 6045 2204
rect 5981 2144 6045 2148
rect 6061 2204 6125 2208
rect 6061 2148 6065 2204
rect 6065 2148 6121 2204
rect 6121 2148 6125 2204
rect 6061 2144 6125 2148
rect 8627 2204 8691 2208
rect 8627 2148 8631 2204
rect 8631 2148 8687 2204
rect 8687 2148 8691 2204
rect 8627 2144 8691 2148
rect 8707 2204 8771 2208
rect 8707 2148 8711 2204
rect 8711 2148 8767 2204
rect 8767 2148 8771 2204
rect 8707 2144 8771 2148
rect 8787 2204 8851 2208
rect 8787 2148 8791 2204
rect 8791 2148 8847 2204
rect 8847 2148 8851 2204
rect 8787 2144 8851 2148
rect 8867 2204 8931 2208
rect 8867 2148 8871 2204
rect 8871 2148 8927 2204
rect 8927 2148 8931 2204
rect 8867 2144 8931 2148
rect 11433 2204 11497 2208
rect 11433 2148 11437 2204
rect 11437 2148 11493 2204
rect 11493 2148 11497 2204
rect 11433 2144 11497 2148
rect 11513 2204 11577 2208
rect 11513 2148 11517 2204
rect 11517 2148 11573 2204
rect 11573 2148 11577 2204
rect 11513 2144 11577 2148
rect 11593 2204 11657 2208
rect 11593 2148 11597 2204
rect 11597 2148 11653 2204
rect 11653 2148 11657 2204
rect 11593 2144 11657 2148
rect 11673 2204 11737 2208
rect 11673 2148 11677 2204
rect 11677 2148 11733 2204
rect 11733 2148 11737 2204
rect 11673 2144 11737 2148
<< metal4 >>
rect 2347 12544 2667 13104
rect 2347 12480 2355 12544
rect 2419 12480 2435 12544
rect 2499 12480 2515 12544
rect 2579 12480 2595 12544
rect 2659 12480 2667 12544
rect 2347 11814 2667 12480
rect 2347 11578 2389 11814
rect 2625 11578 2667 11814
rect 2347 11456 2667 11578
rect 2347 11392 2355 11456
rect 2419 11392 2435 11456
rect 2499 11392 2515 11456
rect 2579 11392 2595 11456
rect 2659 11392 2667 11456
rect 2347 10368 2667 11392
rect 2347 10304 2355 10368
rect 2419 10304 2435 10368
rect 2499 10304 2515 10368
rect 2579 10304 2595 10368
rect 2659 10304 2667 10368
rect 2347 9280 2667 10304
rect 2347 9216 2355 9280
rect 2419 9216 2435 9280
rect 2499 9216 2515 9280
rect 2579 9216 2595 9280
rect 2659 9216 2667 9280
rect 2347 9094 2667 9216
rect 2347 8858 2389 9094
rect 2625 8858 2667 9094
rect 2347 8192 2667 8858
rect 2347 8128 2355 8192
rect 2419 8128 2435 8192
rect 2499 8128 2515 8192
rect 2579 8128 2595 8192
rect 2659 8128 2667 8192
rect 2347 7104 2667 8128
rect 2347 7040 2355 7104
rect 2419 7040 2435 7104
rect 2499 7040 2515 7104
rect 2579 7040 2595 7104
rect 2659 7040 2667 7104
rect 2347 6374 2667 7040
rect 2347 6138 2389 6374
rect 2625 6138 2667 6374
rect 2347 6016 2667 6138
rect 2347 5952 2355 6016
rect 2419 5952 2435 6016
rect 2499 5952 2515 6016
rect 2579 5952 2595 6016
rect 2659 5952 2667 6016
rect 2347 4928 2667 5952
rect 2347 4864 2355 4928
rect 2419 4864 2435 4928
rect 2499 4864 2515 4928
rect 2579 4864 2595 4928
rect 2659 4864 2667 4928
rect 2347 3840 2667 4864
rect 2347 3776 2355 3840
rect 2419 3776 2435 3840
rect 2499 3776 2515 3840
rect 2579 3776 2595 3840
rect 2659 3776 2667 3840
rect 2347 3654 2667 3776
rect 2347 3418 2389 3654
rect 2625 3418 2667 3654
rect 2347 2752 2667 3418
rect 2347 2688 2355 2752
rect 2419 2688 2435 2752
rect 2499 2688 2515 2752
rect 2579 2688 2595 2752
rect 2659 2688 2667 2752
rect 2347 2128 2667 2688
rect 3007 13088 3327 13104
rect 3007 13024 3015 13088
rect 3079 13024 3095 13088
rect 3159 13024 3175 13088
rect 3239 13024 3255 13088
rect 3319 13024 3327 13088
rect 3007 12474 3327 13024
rect 3007 12238 3049 12474
rect 3285 12238 3327 12474
rect 3007 12000 3327 12238
rect 3007 11936 3015 12000
rect 3079 11936 3095 12000
rect 3159 11936 3175 12000
rect 3239 11936 3255 12000
rect 3319 11936 3327 12000
rect 3007 10912 3327 11936
rect 5153 12544 5473 13104
rect 5153 12480 5161 12544
rect 5225 12480 5241 12544
rect 5305 12480 5321 12544
rect 5385 12480 5401 12544
rect 5465 12480 5473 12544
rect 5153 11814 5473 12480
rect 4107 11660 4173 11661
rect 4107 11596 4108 11660
rect 4172 11596 4173 11660
rect 4107 11595 4173 11596
rect 3007 10848 3015 10912
rect 3079 10848 3095 10912
rect 3159 10848 3175 10912
rect 3239 10848 3255 10912
rect 3319 10848 3327 10912
rect 3007 9824 3327 10848
rect 3007 9760 3015 9824
rect 3079 9760 3095 9824
rect 3159 9760 3175 9824
rect 3239 9760 3255 9824
rect 3319 9760 3327 9824
rect 3007 9754 3327 9760
rect 3007 9518 3049 9754
rect 3285 9518 3327 9754
rect 3007 8736 3327 9518
rect 3007 8672 3015 8736
rect 3079 8672 3095 8736
rect 3159 8672 3175 8736
rect 3239 8672 3255 8736
rect 3319 8672 3327 8736
rect 3007 7648 3327 8672
rect 4110 8261 4170 11595
rect 5153 11578 5195 11814
rect 5431 11578 5473 11814
rect 5153 11456 5473 11578
rect 5153 11392 5161 11456
rect 5225 11392 5241 11456
rect 5305 11392 5321 11456
rect 5385 11392 5401 11456
rect 5465 11392 5473 11456
rect 5153 10368 5473 11392
rect 5153 10304 5161 10368
rect 5225 10304 5241 10368
rect 5305 10304 5321 10368
rect 5385 10304 5401 10368
rect 5465 10304 5473 10368
rect 5153 9280 5473 10304
rect 5153 9216 5161 9280
rect 5225 9216 5241 9280
rect 5305 9216 5321 9280
rect 5385 9216 5401 9280
rect 5465 9216 5473 9280
rect 5153 9094 5473 9216
rect 5153 8858 5195 9094
rect 5431 8858 5473 9094
rect 4107 8260 4173 8261
rect 4107 8196 4108 8260
rect 4172 8196 4173 8260
rect 4107 8195 4173 8196
rect 3007 7584 3015 7648
rect 3079 7584 3095 7648
rect 3159 7584 3175 7648
rect 3239 7584 3255 7648
rect 3319 7584 3327 7648
rect 3007 7034 3327 7584
rect 3007 6798 3049 7034
rect 3285 6798 3327 7034
rect 3007 6560 3327 6798
rect 3007 6496 3015 6560
rect 3079 6496 3095 6560
rect 3159 6496 3175 6560
rect 3239 6496 3255 6560
rect 3319 6496 3327 6560
rect 3007 5472 3327 6496
rect 3007 5408 3015 5472
rect 3079 5408 3095 5472
rect 3159 5408 3175 5472
rect 3239 5408 3255 5472
rect 3319 5408 3327 5472
rect 3007 4384 3327 5408
rect 3007 4320 3015 4384
rect 3079 4320 3095 4384
rect 3159 4320 3175 4384
rect 3239 4320 3255 4384
rect 3319 4320 3327 4384
rect 3007 4314 3327 4320
rect 3007 4078 3049 4314
rect 3285 4078 3327 4314
rect 3007 3296 3327 4078
rect 3007 3232 3015 3296
rect 3079 3232 3095 3296
rect 3159 3232 3175 3296
rect 3239 3232 3255 3296
rect 3319 3232 3327 3296
rect 3007 2208 3327 3232
rect 3007 2144 3015 2208
rect 3079 2144 3095 2208
rect 3159 2144 3175 2208
rect 3239 2144 3255 2208
rect 3319 2144 3327 2208
rect 3007 2128 3327 2144
rect 5153 8192 5473 8858
rect 5153 8128 5161 8192
rect 5225 8128 5241 8192
rect 5305 8128 5321 8192
rect 5385 8128 5401 8192
rect 5465 8128 5473 8192
rect 5153 7104 5473 8128
rect 5153 7040 5161 7104
rect 5225 7040 5241 7104
rect 5305 7040 5321 7104
rect 5385 7040 5401 7104
rect 5465 7040 5473 7104
rect 5153 6374 5473 7040
rect 5153 6138 5195 6374
rect 5431 6138 5473 6374
rect 5153 6016 5473 6138
rect 5153 5952 5161 6016
rect 5225 5952 5241 6016
rect 5305 5952 5321 6016
rect 5385 5952 5401 6016
rect 5465 5952 5473 6016
rect 5153 4928 5473 5952
rect 5153 4864 5161 4928
rect 5225 4864 5241 4928
rect 5305 4864 5321 4928
rect 5385 4864 5401 4928
rect 5465 4864 5473 4928
rect 5153 3840 5473 4864
rect 5153 3776 5161 3840
rect 5225 3776 5241 3840
rect 5305 3776 5321 3840
rect 5385 3776 5401 3840
rect 5465 3776 5473 3840
rect 5153 3654 5473 3776
rect 5153 3418 5195 3654
rect 5431 3418 5473 3654
rect 5153 2752 5473 3418
rect 5153 2688 5161 2752
rect 5225 2688 5241 2752
rect 5305 2688 5321 2752
rect 5385 2688 5401 2752
rect 5465 2688 5473 2752
rect 5153 2128 5473 2688
rect 5813 13088 6133 13104
rect 5813 13024 5821 13088
rect 5885 13024 5901 13088
rect 5965 13024 5981 13088
rect 6045 13024 6061 13088
rect 6125 13024 6133 13088
rect 5813 12474 6133 13024
rect 5813 12238 5855 12474
rect 6091 12238 6133 12474
rect 5813 12000 6133 12238
rect 5813 11936 5821 12000
rect 5885 11936 5901 12000
rect 5965 11936 5981 12000
rect 6045 11936 6061 12000
rect 6125 11936 6133 12000
rect 5813 10912 6133 11936
rect 5813 10848 5821 10912
rect 5885 10848 5901 10912
rect 5965 10848 5981 10912
rect 6045 10848 6061 10912
rect 6125 10848 6133 10912
rect 5813 9824 6133 10848
rect 5813 9760 5821 9824
rect 5885 9760 5901 9824
rect 5965 9760 5981 9824
rect 6045 9760 6061 9824
rect 6125 9760 6133 9824
rect 5813 9754 6133 9760
rect 5813 9518 5855 9754
rect 6091 9518 6133 9754
rect 5813 8736 6133 9518
rect 5813 8672 5821 8736
rect 5885 8672 5901 8736
rect 5965 8672 5981 8736
rect 6045 8672 6061 8736
rect 6125 8672 6133 8736
rect 5813 7648 6133 8672
rect 5813 7584 5821 7648
rect 5885 7584 5901 7648
rect 5965 7584 5981 7648
rect 6045 7584 6061 7648
rect 6125 7584 6133 7648
rect 5813 7034 6133 7584
rect 5813 6798 5855 7034
rect 6091 6798 6133 7034
rect 5813 6560 6133 6798
rect 5813 6496 5821 6560
rect 5885 6496 5901 6560
rect 5965 6496 5981 6560
rect 6045 6496 6061 6560
rect 6125 6496 6133 6560
rect 5813 5472 6133 6496
rect 5813 5408 5821 5472
rect 5885 5408 5901 5472
rect 5965 5408 5981 5472
rect 6045 5408 6061 5472
rect 6125 5408 6133 5472
rect 5813 4384 6133 5408
rect 5813 4320 5821 4384
rect 5885 4320 5901 4384
rect 5965 4320 5981 4384
rect 6045 4320 6061 4384
rect 6125 4320 6133 4384
rect 5813 4314 6133 4320
rect 5813 4078 5855 4314
rect 6091 4078 6133 4314
rect 5813 3296 6133 4078
rect 5813 3232 5821 3296
rect 5885 3232 5901 3296
rect 5965 3232 5981 3296
rect 6045 3232 6061 3296
rect 6125 3232 6133 3296
rect 5813 2208 6133 3232
rect 5813 2144 5821 2208
rect 5885 2144 5901 2208
rect 5965 2144 5981 2208
rect 6045 2144 6061 2208
rect 6125 2144 6133 2208
rect 5813 2128 6133 2144
rect 7959 12544 8279 13104
rect 7959 12480 7967 12544
rect 8031 12480 8047 12544
rect 8111 12480 8127 12544
rect 8191 12480 8207 12544
rect 8271 12480 8279 12544
rect 7959 11814 8279 12480
rect 7959 11578 8001 11814
rect 8237 11578 8279 11814
rect 7959 11456 8279 11578
rect 7959 11392 7967 11456
rect 8031 11392 8047 11456
rect 8111 11392 8127 11456
rect 8191 11392 8207 11456
rect 8271 11392 8279 11456
rect 7959 10368 8279 11392
rect 7959 10304 7967 10368
rect 8031 10304 8047 10368
rect 8111 10304 8127 10368
rect 8191 10304 8207 10368
rect 8271 10304 8279 10368
rect 7959 9280 8279 10304
rect 7959 9216 7967 9280
rect 8031 9216 8047 9280
rect 8111 9216 8127 9280
rect 8191 9216 8207 9280
rect 8271 9216 8279 9280
rect 7959 9094 8279 9216
rect 7959 8858 8001 9094
rect 8237 8858 8279 9094
rect 7959 8192 8279 8858
rect 7959 8128 7967 8192
rect 8031 8128 8047 8192
rect 8111 8128 8127 8192
rect 8191 8128 8207 8192
rect 8271 8128 8279 8192
rect 7959 7104 8279 8128
rect 7959 7040 7967 7104
rect 8031 7040 8047 7104
rect 8111 7040 8127 7104
rect 8191 7040 8207 7104
rect 8271 7040 8279 7104
rect 7959 6374 8279 7040
rect 7959 6138 8001 6374
rect 8237 6138 8279 6374
rect 7959 6016 8279 6138
rect 7959 5952 7967 6016
rect 8031 5952 8047 6016
rect 8111 5952 8127 6016
rect 8191 5952 8207 6016
rect 8271 5952 8279 6016
rect 7959 4928 8279 5952
rect 7959 4864 7967 4928
rect 8031 4864 8047 4928
rect 8111 4864 8127 4928
rect 8191 4864 8207 4928
rect 8271 4864 8279 4928
rect 7959 3840 8279 4864
rect 7959 3776 7967 3840
rect 8031 3776 8047 3840
rect 8111 3776 8127 3840
rect 8191 3776 8207 3840
rect 8271 3776 8279 3840
rect 7959 3654 8279 3776
rect 7959 3418 8001 3654
rect 8237 3418 8279 3654
rect 7959 2752 8279 3418
rect 7959 2688 7967 2752
rect 8031 2688 8047 2752
rect 8111 2688 8127 2752
rect 8191 2688 8207 2752
rect 8271 2688 8279 2752
rect 7959 2128 8279 2688
rect 8619 13088 8939 13104
rect 8619 13024 8627 13088
rect 8691 13024 8707 13088
rect 8771 13024 8787 13088
rect 8851 13024 8867 13088
rect 8931 13024 8939 13088
rect 8619 12474 8939 13024
rect 8619 12238 8661 12474
rect 8897 12238 8939 12474
rect 8619 12000 8939 12238
rect 8619 11936 8627 12000
rect 8691 11936 8707 12000
rect 8771 11936 8787 12000
rect 8851 11936 8867 12000
rect 8931 11936 8939 12000
rect 8619 10912 8939 11936
rect 8619 10848 8627 10912
rect 8691 10848 8707 10912
rect 8771 10848 8787 10912
rect 8851 10848 8867 10912
rect 8931 10848 8939 10912
rect 8619 9824 8939 10848
rect 8619 9760 8627 9824
rect 8691 9760 8707 9824
rect 8771 9760 8787 9824
rect 8851 9760 8867 9824
rect 8931 9760 8939 9824
rect 8619 9754 8939 9760
rect 8619 9518 8661 9754
rect 8897 9518 8939 9754
rect 8619 8736 8939 9518
rect 8619 8672 8627 8736
rect 8691 8672 8707 8736
rect 8771 8672 8787 8736
rect 8851 8672 8867 8736
rect 8931 8672 8939 8736
rect 8619 7648 8939 8672
rect 8619 7584 8627 7648
rect 8691 7584 8707 7648
rect 8771 7584 8787 7648
rect 8851 7584 8867 7648
rect 8931 7584 8939 7648
rect 8619 7034 8939 7584
rect 8619 6798 8661 7034
rect 8897 6798 8939 7034
rect 8619 6560 8939 6798
rect 8619 6496 8627 6560
rect 8691 6496 8707 6560
rect 8771 6496 8787 6560
rect 8851 6496 8867 6560
rect 8931 6496 8939 6560
rect 8619 5472 8939 6496
rect 8619 5408 8627 5472
rect 8691 5408 8707 5472
rect 8771 5408 8787 5472
rect 8851 5408 8867 5472
rect 8931 5408 8939 5472
rect 8619 4384 8939 5408
rect 8619 4320 8627 4384
rect 8691 4320 8707 4384
rect 8771 4320 8787 4384
rect 8851 4320 8867 4384
rect 8931 4320 8939 4384
rect 8619 4314 8939 4320
rect 8619 4078 8661 4314
rect 8897 4078 8939 4314
rect 8619 3296 8939 4078
rect 8619 3232 8627 3296
rect 8691 3232 8707 3296
rect 8771 3232 8787 3296
rect 8851 3232 8867 3296
rect 8931 3232 8939 3296
rect 8619 2208 8939 3232
rect 8619 2144 8627 2208
rect 8691 2144 8707 2208
rect 8771 2144 8787 2208
rect 8851 2144 8867 2208
rect 8931 2144 8939 2208
rect 8619 2128 8939 2144
rect 10765 12544 11085 13104
rect 10765 12480 10773 12544
rect 10837 12480 10853 12544
rect 10917 12480 10933 12544
rect 10997 12480 11013 12544
rect 11077 12480 11085 12544
rect 10765 11814 11085 12480
rect 10765 11578 10807 11814
rect 11043 11578 11085 11814
rect 10765 11456 11085 11578
rect 10765 11392 10773 11456
rect 10837 11392 10853 11456
rect 10917 11392 10933 11456
rect 10997 11392 11013 11456
rect 11077 11392 11085 11456
rect 10765 10368 11085 11392
rect 10765 10304 10773 10368
rect 10837 10304 10853 10368
rect 10917 10304 10933 10368
rect 10997 10304 11013 10368
rect 11077 10304 11085 10368
rect 10765 9280 11085 10304
rect 10765 9216 10773 9280
rect 10837 9216 10853 9280
rect 10917 9216 10933 9280
rect 10997 9216 11013 9280
rect 11077 9216 11085 9280
rect 10765 9094 11085 9216
rect 10765 8858 10807 9094
rect 11043 8858 11085 9094
rect 10765 8192 11085 8858
rect 10765 8128 10773 8192
rect 10837 8128 10853 8192
rect 10917 8128 10933 8192
rect 10997 8128 11013 8192
rect 11077 8128 11085 8192
rect 10765 7104 11085 8128
rect 10765 7040 10773 7104
rect 10837 7040 10853 7104
rect 10917 7040 10933 7104
rect 10997 7040 11013 7104
rect 11077 7040 11085 7104
rect 10765 6374 11085 7040
rect 10765 6138 10807 6374
rect 11043 6138 11085 6374
rect 10765 6016 11085 6138
rect 10765 5952 10773 6016
rect 10837 5952 10853 6016
rect 10917 5952 10933 6016
rect 10997 5952 11013 6016
rect 11077 5952 11085 6016
rect 10765 4928 11085 5952
rect 10765 4864 10773 4928
rect 10837 4864 10853 4928
rect 10917 4864 10933 4928
rect 10997 4864 11013 4928
rect 11077 4864 11085 4928
rect 10765 3840 11085 4864
rect 10765 3776 10773 3840
rect 10837 3776 10853 3840
rect 10917 3776 10933 3840
rect 10997 3776 11013 3840
rect 11077 3776 11085 3840
rect 10765 3654 11085 3776
rect 10765 3418 10807 3654
rect 11043 3418 11085 3654
rect 10765 2752 11085 3418
rect 10765 2688 10773 2752
rect 10837 2688 10853 2752
rect 10917 2688 10933 2752
rect 10997 2688 11013 2752
rect 11077 2688 11085 2752
rect 10765 2128 11085 2688
rect 11425 13088 11745 13104
rect 11425 13024 11433 13088
rect 11497 13024 11513 13088
rect 11577 13024 11593 13088
rect 11657 13024 11673 13088
rect 11737 13024 11745 13088
rect 11425 12474 11745 13024
rect 11425 12238 11467 12474
rect 11703 12238 11745 12474
rect 11425 12000 11745 12238
rect 11425 11936 11433 12000
rect 11497 11936 11513 12000
rect 11577 11936 11593 12000
rect 11657 11936 11673 12000
rect 11737 11936 11745 12000
rect 11425 10912 11745 11936
rect 11425 10848 11433 10912
rect 11497 10848 11513 10912
rect 11577 10848 11593 10912
rect 11657 10848 11673 10912
rect 11737 10848 11745 10912
rect 11425 9824 11745 10848
rect 11425 9760 11433 9824
rect 11497 9760 11513 9824
rect 11577 9760 11593 9824
rect 11657 9760 11673 9824
rect 11737 9760 11745 9824
rect 11425 9754 11745 9760
rect 11425 9518 11467 9754
rect 11703 9518 11745 9754
rect 11425 8736 11745 9518
rect 11425 8672 11433 8736
rect 11497 8672 11513 8736
rect 11577 8672 11593 8736
rect 11657 8672 11673 8736
rect 11737 8672 11745 8736
rect 11425 7648 11745 8672
rect 11425 7584 11433 7648
rect 11497 7584 11513 7648
rect 11577 7584 11593 7648
rect 11657 7584 11673 7648
rect 11737 7584 11745 7648
rect 11425 7034 11745 7584
rect 11425 6798 11467 7034
rect 11703 6798 11745 7034
rect 11425 6560 11745 6798
rect 11425 6496 11433 6560
rect 11497 6496 11513 6560
rect 11577 6496 11593 6560
rect 11657 6496 11673 6560
rect 11737 6496 11745 6560
rect 11425 5472 11745 6496
rect 11425 5408 11433 5472
rect 11497 5408 11513 5472
rect 11577 5408 11593 5472
rect 11657 5408 11673 5472
rect 11737 5408 11745 5472
rect 11425 4384 11745 5408
rect 11425 4320 11433 4384
rect 11497 4320 11513 4384
rect 11577 4320 11593 4384
rect 11657 4320 11673 4384
rect 11737 4320 11745 4384
rect 11425 4314 11745 4320
rect 11425 4078 11467 4314
rect 11703 4078 11745 4314
rect 11425 3296 11745 4078
rect 11425 3232 11433 3296
rect 11497 3232 11513 3296
rect 11577 3232 11593 3296
rect 11657 3232 11673 3296
rect 11737 3232 11745 3296
rect 11425 2208 11745 3232
rect 11425 2144 11433 2208
rect 11497 2144 11513 2208
rect 11577 2144 11593 2208
rect 11657 2144 11673 2208
rect 11737 2144 11745 2208
rect 11425 2128 11745 2144
<< via4 >>
rect 2389 11578 2625 11814
rect 2389 8858 2625 9094
rect 2389 6138 2625 6374
rect 2389 3418 2625 3654
rect 3049 12238 3285 12474
rect 3049 9518 3285 9754
rect 5195 11578 5431 11814
rect 5195 8858 5431 9094
rect 3049 6798 3285 7034
rect 3049 4078 3285 4314
rect 5195 6138 5431 6374
rect 5195 3418 5431 3654
rect 5855 12238 6091 12474
rect 5855 9518 6091 9754
rect 5855 6798 6091 7034
rect 5855 4078 6091 4314
rect 8001 11578 8237 11814
rect 8001 8858 8237 9094
rect 8001 6138 8237 6374
rect 8001 3418 8237 3654
rect 8661 12238 8897 12474
rect 8661 9518 8897 9754
rect 8661 6798 8897 7034
rect 8661 4078 8897 4314
rect 10807 11578 11043 11814
rect 10807 8858 11043 9094
rect 10807 6138 11043 6374
rect 10807 3418 11043 3654
rect 11467 12238 11703 12474
rect 11467 9518 11703 9754
rect 11467 6798 11703 7034
rect 11467 4078 11703 4314
<< metal5 >>
rect 1056 12474 12376 12516
rect 1056 12238 3049 12474
rect 3285 12238 5855 12474
rect 6091 12238 8661 12474
rect 8897 12238 11467 12474
rect 11703 12238 12376 12474
rect 1056 12196 12376 12238
rect 1056 11814 12376 11856
rect 1056 11578 2389 11814
rect 2625 11578 5195 11814
rect 5431 11578 8001 11814
rect 8237 11578 10807 11814
rect 11043 11578 12376 11814
rect 1056 11536 12376 11578
rect 1056 9754 12376 9796
rect 1056 9518 3049 9754
rect 3285 9518 5855 9754
rect 6091 9518 8661 9754
rect 8897 9518 11467 9754
rect 11703 9518 12376 9754
rect 1056 9476 12376 9518
rect 1056 9094 12376 9136
rect 1056 8858 2389 9094
rect 2625 8858 5195 9094
rect 5431 8858 8001 9094
rect 8237 8858 10807 9094
rect 11043 8858 12376 9094
rect 1056 8816 12376 8858
rect 1056 7034 12376 7076
rect 1056 6798 3049 7034
rect 3285 6798 5855 7034
rect 6091 6798 8661 7034
rect 8897 6798 11467 7034
rect 11703 6798 12376 7034
rect 1056 6756 12376 6798
rect 1056 6374 12376 6416
rect 1056 6138 2389 6374
rect 2625 6138 5195 6374
rect 5431 6138 8001 6374
rect 8237 6138 10807 6374
rect 11043 6138 12376 6374
rect 1056 6096 12376 6138
rect 1056 4314 12376 4356
rect 1056 4078 3049 4314
rect 3285 4078 5855 4314
rect 6091 4078 8661 4314
rect 8897 4078 11467 4314
rect 11703 4078 12376 4314
rect 1056 4036 12376 4078
rect 1056 3654 12376 3696
rect 1056 3418 2389 3654
rect 2625 3418 5195 3654
rect 5431 3418 8001 3654
rect 8237 3418 10807 3654
rect 11043 3418 12376 3654
rect 1056 3376 12376 3418
use sky130_fd_sc_hd__dlymetal6s2s_1  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8740 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1704896540
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _124_
timestamp 1704896540
transform 1 0 8464 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _125_
timestamp 1704896540
transform 1 0 8280 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _127_
timestamp 1704896540
transform 1 0 8740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9752 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1704896540
transform -1 0 5428 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _131_
timestamp 1704896540
transform -1 0 8464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9936 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9936 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1704896540
transform 1 0 10120 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11316 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _136_
timestamp 1704896540
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _137_
timestamp 1704896540
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10580 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10396 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _141_
timestamp 1704896540
transform -1 0 10948 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11960 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _146_
timestamp 1704896540
transform 1 0 11316 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _147_
timestamp 1704896540
transform -1 0 12052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_2  _148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9752 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _150_
timestamp 1704896540
transform 1 0 9844 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9292 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a311oi_2  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11132 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _154_
timestamp 1704896540
transform 1 0 7176 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _156_
timestamp 1704896540
transform -1 0 8280 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _157_
timestamp 1704896540
transform -1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1704896540
transform -1 0 7360 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _160_
timestamp 1704896540
transform -1 0 6256 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1704896540
transform 1 0 3864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o311ai_2  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5060 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1704896540
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _164_
timestamp 1704896540
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _165_
timestamp 1704896540
transform -1 0 6164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _166_
timestamp 1704896540
transform 1 0 5428 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _167_
timestamp 1704896540
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7820 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _169_
timestamp 1704896540
transform 1 0 4508 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1704896540
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _171_
timestamp 1704896540
transform 1 0 11224 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _172_
timestamp 1704896540
transform -1 0 10764 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _173_
timestamp 1704896540
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _174_
timestamp 1704896540
transform -1 0 5980 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _175_
timestamp 1704896540
transform 1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _176_
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1704896540
transform -1 0 11408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10488 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _182_
timestamp 1704896540
transform -1 0 10488 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _183_
timestamp 1704896540
transform -1 0 6256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _184_
timestamp 1704896540
transform 1 0 4968 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 1704896540
transform -1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5060 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _187_
timestamp 1704896540
transform 1 0 10304 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _188_
timestamp 1704896540
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _189_
timestamp 1704896540
transform 1 0 7084 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _190_
timestamp 1704896540
transform -1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _192_
timestamp 1704896540
transform -1 0 9292 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7728 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _196_
timestamp 1704896540
transform 1 0 9752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _197_
timestamp 1704896540
transform 1 0 9108 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _198_
timestamp 1704896540
transform -1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _199_
timestamp 1704896540
transform -1 0 7084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _200_
timestamp 1704896540
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _201_
timestamp 1704896540
transform 1 0 7636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _202_
timestamp 1704896540
transform 1 0 9568 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _204_
timestamp 1704896540
transform -1 0 6532 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a311o_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _206_
timestamp 1704896540
transform 1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _207_
timestamp 1704896540
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1704896540
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _209_
timestamp 1704896540
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _210_
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _211_
timestamp 1704896540
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7268 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _213_
timestamp 1704896540
transform 1 0 5520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _214_
timestamp 1704896540
transform -1 0 6256 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _215_
timestamp 1704896540
transform 1 0 6256 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _216_
timestamp 1704896540
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _218_
timestamp 1704896540
transform -1 0 10396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _219_
timestamp 1704896540
transform -1 0 8464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _220_
timestamp 1704896540
transform -1 0 9660 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _222_
timestamp 1704896540
transform 1 0 3680 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1704896540
transform 1 0 2300 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1704896540
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1704896540
transform 1 0 2300 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1704896540
transform 1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1704896540
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1704896540
transform -1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1704896540
transform 1 0 5060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1704896540
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1704896540
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1704896540
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1704896540
transform -1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1704896540
transform -1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1704896540
transform 1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1704896540
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3404 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 1704896540
transform 1 0 1840 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _243_
timestamp 1704896540
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 1704896540
transform 1 0 6992 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _246_
timestamp 1704896540
transform 1 0 6992 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _247_
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _248_
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 1704896540
transform 1 0 2576 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _250_
timestamp 1704896540
transform -1 0 3680 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 5612 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform -1 0 5060 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinvlp_2  clkload0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1704896540
transform -1 0 5520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1704896540
transform -1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1704896540
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_70
timestamp 1704896540
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_30
timestamp 1704896540
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1704896540
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_84 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8832 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_92
timestamp 1704896540
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_97
timestamp 1704896540
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_33
timestamp 1704896540
transform 1 0 4140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_45
timestamp 1704896540
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_63
timestamp 1704896540
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_77
timestamp 1704896540
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_105
timestamp 1704896540
transform 1 0 10764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_113
timestamp 1704896540
transform 1 0 11500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_11
timestamp 1704896540
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_22
timestamp 1704896540
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_26
timestamp 1704896540
transform 1 0 3496 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_37
timestamp 1704896540
transform 1 0 4508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_45
timestamp 1704896540
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1704896540
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_72
timestamp 1704896540
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_82
timestamp 1704896540
transform 1 0 8648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_90
timestamp 1704896540
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_98
timestamp 1704896540
transform 1 0 10120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_118
timestamp 1704896540
transform 1 0 11960 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_48
timestamp 1704896540
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_60
timestamp 1704896540
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_72
timestamp 1704896540
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_92
timestamp 1704896540
transform 1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_114
timestamp 1704896540
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_118
timestamp 1704896540
transform 1 0 11960 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_62
timestamp 1704896540
transform 1 0 6808 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_70
timestamp 1704896540
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_76
timestamp 1704896540
transform 1 0 8096 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_88
timestamp 1704896540
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_100
timestamp 1704896540
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_59
timestamp 1704896540
transform 1 0 6532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_63
timestamp 1704896540
transform 1 0 6900 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_97
timestamp 1704896540
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_106
timestamp 1704896540
transform 1 0 10856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_114
timestamp 1704896540
transform 1 0 11592 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_7
timestamp 1704896540
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_35
timestamp 1704896540
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_47
timestamp 1704896540
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_77
timestamp 1704896540
transform 1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_83
timestamp 1704896540
transform 1 0 8740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_95
timestamp 1704896540
transform 1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_11
timestamp 1704896540
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_33
timestamp 1704896540
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_62
timestamp 1704896540
transform 1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_70
timestamp 1704896540
transform 1 0 7544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 1704896540
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_98
timestamp 1704896540
transform 1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_118
timestamp 1704896540
transform 1 0 11960 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_36
timestamp 1704896540
transform 1 0 4416 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_42
timestamp 1704896540
transform 1 0 4968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_70
timestamp 1704896540
transform 1 0 7544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_74
timestamp 1704896540
transform 1 0 7912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 1704896540
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_7
timestamp 1704896540
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_13
timestamp 1704896540
transform 1 0 2300 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_32
timestamp 1704896540
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_54
timestamp 1704896540
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_64
timestamp 1704896540
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_76
timestamp 1704896540
transform 1 0 8096 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1704896540
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_103
timestamp 1704896540
transform 1 0 10580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_115
timestamp 1704896540
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_25
timestamp 1704896540
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_37
timestamp 1704896540
transform 1 0 4508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_66
timestamp 1704896540
transform 1 0 7176 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_78
timestamp 1704896540
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_89
timestamp 1704896540
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_101
timestamp 1704896540
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1704896540
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_11
timestamp 1704896540
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_17
timestamp 1704896540
transform 1 0 2668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_21
timestamp 1704896540
transform 1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_54
timestamp 1704896540
transform 1 0 6072 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_66
timestamp 1704896540
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1704896540
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_88
timestamp 1704896540
transform 1 0 9200 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_103
timestamp 1704896540
transform 1 0 10580 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_43
timestamp 1704896540
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 1704896540
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_68
timestamp 1704896540
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_80
timestamp 1704896540
transform 1 0 8464 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_96
timestamp 1704896540
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_108
timestamp 1704896540
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_7
timestamp 1704896540
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1704896540
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_56
timestamp 1704896540
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_68
timestamp 1704896540
transform 1 0 7360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_76
timestamp 1704896540
transform 1 0 8096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_80
timestamp 1704896540
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_99
timestamp 1704896540
transform 1 0 10212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_111
timestamp 1704896540
transform 1 0 11316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_115
timestamp 1704896540
transform 1 0 11684 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_26
timestamp 1704896540
transform 1 0 3496 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_34
timestamp 1704896540
transform 1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1704896540
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_63
timestamp 1704896540
transform 1 0 6900 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_71
timestamp 1704896540
transform 1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_85
timestamp 1704896540
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_97
timestamp 1704896540
transform 1 0 10028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_7
timestamp 1704896540
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_19
timestamp 1704896540
transform 1 0 2852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 1704896540
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_48
timestamp 1704896540
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_65
timestamp 1704896540
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_69
timestamp 1704896540
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_74
timestamp 1704896540
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1704896540
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_117
timestamp 1704896540
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_11
timestamp 1704896540
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_36
timestamp 1704896540
transform 1 0 4416 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_45
timestamp 1704896540
transform 1 0 5244 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1704896540
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_65
timestamp 1704896540
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_86
timestamp 1704896540
transform 1 0 9016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1704896540
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_48
timestamp 1704896540
transform 1 0 5520 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_61
timestamp 1704896540
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_65
timestamp 1704896540
transform 1 0 7084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 1704896540
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_93
timestamp 1704896540
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_105
timestamp 1704896540
transform 1 0 10764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_117
timestamp 1704896540
transform 1 0 11868 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3588 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_29
timestamp 1704896540
transform 1 0 3772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_41
timestamp 1704896540
transform 1 0 4876 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_49
timestamp 1704896540
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1704896540
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_69
timestamp 1704896540
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_76
timestamp 1704896540
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_83
timestamp 1704896540
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_85
timestamp 1704896540
transform 1 0 8924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_97
timestamp 1704896540
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1704896540
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 2392 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1704896540
transform -1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 11776 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform -1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1704896540
transform 1 0 8464 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1704896540
transform -1 0 8096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1704896540
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1704896540
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1704896540
transform -1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1704896540
transform -1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1704896540
transform 1 0 11684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1704896540
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1704896540
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1704896540
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_20
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_21
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_22
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_23
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_24
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 12328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_25
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_26
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_27
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_28
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_29
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_30
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_31
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_32
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_33
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 12328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_34
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_35
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 12328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_36
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_37
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 12328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_38
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 12328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_39
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 12328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_41
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_42
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_43
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_50
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_51
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_52
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_53
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_54
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_56
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_57
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_58
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_59
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_60
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_61
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_62
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_63
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_64
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_65
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_66
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_67
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_68
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_69
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_70
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_71
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_72
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_73
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_74
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_75
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_76
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_77
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_78
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_79
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_80
timestamp 1704896540
transform 1 0 3680 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_81
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_82
timestamp 1704896540
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_83
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
<< labels >>
flabel metal4 s 3007 2128 3327 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5813 2128 6133 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8619 2128 8939 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11425 2128 11745 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4036 12376 4356 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6756 12376 7076 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9476 12376 9796 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 12196 12376 12516 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2347 2128 2667 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5153 2128 5473 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7959 2128 8279 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10765 2128 11085 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3376 12376 3696 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 6096 12376 6416 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8816 12376 9136 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 11536 12376 11856 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 current[0]
port 3 nsew signal input
flabel metal3 s 12699 3408 13499 3528 0 FreeSans 480 0 0 0 current[1]
port 4 nsew signal input
flabel metal3 s 12699 4768 13499 4888 0 FreeSans 480 0 0 0 current[2]
port 5 nsew signal input
flabel metal3 s 12699 5448 13499 5568 0 FreeSans 480 0 0 0 current[3]
port 6 nsew signal input
flabel metal3 s 12699 9528 13499 9648 0 FreeSans 480 0 0 0 current[4]
port 7 nsew signal input
flabel metal2 s 8390 14843 8446 15643 0 FreeSans 224 90 0 0 current[5]
port 8 nsew signal input
flabel metal2 s 7746 14843 7802 15643 0 FreeSans 224 90 0 0 current[6]
port 9 nsew signal input
flabel metal2 s 7102 14843 7158 15643 0 FreeSans 224 90 0 0 current[7]
port 10 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 reset
port 11 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 spike
port 12 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 voltage[0]
port 13 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 voltage[1]
port 14 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 voltage[2]
port 15 nsew signal output
flabel metal3 s 12699 6128 13499 6248 0 FreeSans 480 0 0 0 voltage[3]
port 16 nsew signal output
flabel metal3 s 12699 8848 13499 8968 0 FreeSans 480 0 0 0 voltage[4]
port 17 nsew signal output
flabel metal2 s 6458 14843 6514 15643 0 FreeSans 224 90 0 0 voltage[5]
port 18 nsew signal output
flabel metal2 s 5814 14843 5870 15643 0 FreeSans 224 90 0 0 voltage[6]
port 19 nsew signal output
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 voltage[7]
port 20 nsew signal output
rlabel metal1 6716 13056 6716 13056 0 VGND
rlabel metal1 6716 12512 6716 12512 0 VPWR
rlabel metal1 1978 8425 1978 8425 0 _000_
rlabel metal2 3726 3298 3726 3298 0 _001_
rlabel metal1 3917 6358 3917 6358 0 _002_
rlabel metal1 5382 2618 5382 2618 0 _003_
rlabel metal2 8050 3230 8050 3230 0 _004_
rlabel metal2 4646 4998 4646 4998 0 _005_
rlabel metal1 8142 5338 8142 5338 0 _006_
rlabel metal1 2852 9146 2852 9146 0 _007_
rlabel metal1 3135 10710 3135 10710 0 _008_
rlabel metal1 3312 11322 3312 11322 0 _009_
rlabel metal1 2392 11866 2392 11866 0 _010_
rlabel via1 1697 3026 1697 3026 0 _011_
rlabel via1 1697 5678 1697 5678 0 _012_
rlabel metal1 3128 8058 3128 8058 0 _013_
rlabel metal1 4462 3128 4462 3128 0 _014_
rlabel metal2 7314 3230 7314 3230 0 _015_
rlabel metal1 4416 4794 4416 4794 0 _016_
rlabel metal2 7314 6188 7314 6188 0 _017_
rlabel metal1 2070 9146 2070 9146 0 _018_
rlabel metal1 1702 10744 1702 10744 0 _019_
rlabel metal1 3726 11662 3726 11662 0 _020_
rlabel metal2 4554 11730 4554 11730 0 _021_
rlabel metal2 5566 10404 5566 10404 0 _022_
rlabel metal1 6394 10506 6394 10506 0 _023_
rlabel metal2 6394 11254 6394 11254 0 _024_
rlabel metal1 4738 11696 4738 11696 0 _025_
rlabel metal2 10810 10880 10810 10880 0 _026_
rlabel metal2 10442 11016 10442 11016 0 _027_
rlabel metal1 10442 11152 10442 11152 0 _028_
rlabel metal1 5290 11118 5290 11118 0 _029_
rlabel metal1 5474 10064 5474 10064 0 _030_
rlabel metal1 5060 10234 5060 10234 0 _031_
rlabel metal1 5474 11084 5474 11084 0 _032_
rlabel metal2 10350 7412 10350 7412 0 _033_
rlabel metal1 9752 8398 9752 8398 0 _034_
rlabel metal1 7084 7514 7084 7514 0 _035_
rlabel metal2 6854 8262 6854 8262 0 _036_
rlabel metal1 8786 8364 8786 8364 0 _037_
rlabel metal1 8740 8602 8740 8602 0 _038_
rlabel metal1 2622 9010 2622 9010 0 _039_
rlabel metal1 10396 6698 10396 6698 0 _040_
rlabel metal1 8326 7344 8326 7344 0 _041_
rlabel metal1 8786 6970 8786 6970 0 _042_
rlabel metal1 6624 6970 6624 6970 0 _043_
rlabel metal1 8510 7412 8510 7412 0 _044_
rlabel metal2 7866 6970 7866 6970 0 _045_
rlabel metal1 9476 4250 9476 4250 0 _046_
rlabel metal1 5382 4624 5382 4624 0 _047_
rlabel metal1 5566 4590 5566 4590 0 _048_
rlabel metal1 7406 3706 7406 3706 0 _049_
rlabel metal2 7498 3706 7498 3706 0 _050_
rlabel metal1 7682 3638 7682 3638 0 _051_
rlabel metal1 9660 3162 9660 3162 0 _052_
rlabel metal2 8970 3910 8970 3910 0 _053_
rlabel metal2 7590 3740 7590 3740 0 _054_
rlabel metal2 6486 3740 6486 3740 0 _055_
rlabel metal1 6762 3468 6762 3468 0 _056_
rlabel via1 4094 7293 4094 7293 0 _057_
rlabel metal1 9752 4794 9752 4794 0 _058_
rlabel metal2 9614 8942 9614 8942 0 _059_
rlabel metal1 4186 7276 4186 7276 0 _060_
rlabel metal2 2714 5576 2714 5576 0 _061_
rlabel metal2 1794 3706 1794 3706 0 _062_
rlabel metal1 2208 6630 2208 6630 0 _063_
rlabel metal1 4600 2414 4600 2414 0 _064_
rlabel metal2 2806 7242 2806 7242 0 _065_
rlabel metal2 9154 7650 9154 7650 0 _066_
rlabel metal2 6578 10880 6578 10880 0 _067_
rlabel metal1 6578 3638 6578 3638 0 _068_
rlabel metal1 8648 8466 8648 8466 0 _069_
rlabel metal1 9844 11662 9844 11662 0 _070_
rlabel metal1 8050 11866 8050 11866 0 _071_
rlabel metal1 8786 11764 8786 11764 0 _072_
rlabel metal1 9522 11696 9522 11696 0 _073_
rlabel metal2 9338 11968 9338 11968 0 _074_
rlabel metal1 6578 8398 6578 8398 0 _075_
rlabel metal2 6026 10098 6026 10098 0 _076_
rlabel metal2 9338 9758 9338 9758 0 _077_
rlabel metal2 11362 10030 11362 10030 0 _078_
rlabel metal1 10994 8874 10994 8874 0 _079_
rlabel metal1 10764 6358 10764 6358 0 _080_
rlabel metal1 11500 9078 11500 9078 0 _081_
rlabel metal2 11270 6562 11270 6562 0 _082_
rlabel metal1 10856 6290 10856 6290 0 _083_
rlabel metal2 10718 6596 10718 6596 0 _084_
rlabel metal1 11408 4114 11408 4114 0 _085_
rlabel metal2 9982 4046 9982 4046 0 _086_
rlabel metal1 9798 2992 9798 2992 0 _087_
rlabel metal1 9568 3570 9568 3570 0 _088_
rlabel metal1 11178 3502 11178 3502 0 _089_
rlabel metal1 9706 4522 9706 4522 0 _090_
rlabel metal1 11454 6970 11454 6970 0 _091_
rlabel metal1 12006 8908 12006 8908 0 _092_
rlabel metal2 10534 8500 10534 8500 0 _093_
rlabel metal1 10212 7514 10212 7514 0 _094_
rlabel metal2 9890 12002 9890 12002 0 _095_
rlabel metal1 10396 12206 10396 12206 0 _096_
rlabel metal1 10442 10574 10442 10574 0 _097_
rlabel metal1 8234 11560 8234 11560 0 _098_
rlabel metal1 6992 12274 6992 12274 0 _099_
rlabel metal1 8004 11730 8004 11730 0 _100_
rlabel metal1 7590 11322 7590 11322 0 _101_
rlabel metal1 7590 11628 7590 11628 0 _102_
rlabel metal2 8326 6596 8326 6596 0 _103_
rlabel metal1 5704 8330 5704 8330 0 _104_
rlabel metal1 6394 5202 6394 5202 0 _105_
rlabel metal1 5796 5678 5796 5678 0 _106_
rlabel metal1 5750 7446 5750 7446 0 _107_
rlabel metal1 6808 7786 6808 7786 0 _108_
rlabel metal1 6210 4046 6210 4046 0 _109_
rlabel metal2 6394 5474 6394 5474 0 _110_
rlabel metal1 5888 8602 5888 8602 0 _111_
rlabel metal2 5934 9248 5934 9248 0 _112_
rlabel metal2 7314 10642 7314 10642 0 _113_
rlabel metal2 4738 11322 4738 11322 0 _114_
rlabel metal1 5658 11662 5658 11662 0 _115_
rlabel metal2 11270 11764 11270 11764 0 _116_
rlabel metal1 5842 11764 5842 11764 0 _117_
rlabel viali 6210 10031 6210 10031 0 _118_
rlabel metal4 4140 9928 4140 9928 0 clk
rlabel metal1 5290 8058 5290 8058 0 clknet_0_clk
rlabel metal1 2208 6222 2208 6222 0 clknet_1_0__leaf_clk
rlabel metal2 2622 12002 2622 12002 0 clknet_1_1__leaf_clk
rlabel metal2 5842 1027 5842 1027 0 current[0]
rlabel via2 11914 3451 11914 3451 0 current[1]
rlabel metal2 12006 5015 12006 5015 0 current[2]
rlabel metal2 12006 5593 12006 5593 0 current[3]
rlabel metal2 12006 9809 12006 9809 0 current[4]
rlabel metal1 8556 12818 8556 12818 0 current[5]
rlabel metal1 7820 12818 7820 12818 0 current[6]
rlabel metal1 7176 12818 7176 12818 0 current[7]
rlabel metal1 6164 2618 6164 2618 0 net1
rlabel metal1 1656 7854 1656 7854 0 net10
rlabel metal1 8602 3434 8602 3434 0 net11
rlabel metal1 9016 4182 9016 4182 0 net12
rlabel metal1 7774 2482 7774 2482 0 net13
rlabel metal2 8694 6086 8694 6086 0 net14
rlabel metal2 5566 8908 5566 8908 0 net15
rlabel metal1 5198 10642 5198 10642 0 net16
rlabel metal1 5704 12818 5704 12818 0 net17
rlabel metal1 1656 10030 1656 10030 0 net18
rlabel metal1 7866 12172 7866 12172 0 net19
rlabel metal1 10626 4148 10626 4148 0 net2
rlabel metal1 7590 2414 7590 2414 0 net20
rlabel metal2 2898 6052 2898 6052 0 net21
rlabel metal2 2162 3298 2162 3298 0 net22
rlabel metal1 3220 7854 3220 7854 0 net23
rlabel metal2 10718 4794 10718 4794 0 net3
rlabel metal1 10120 6290 10120 6290 0 net4
rlabel metal1 9016 9962 9016 9962 0 net5
rlabel metal1 8234 10676 8234 10676 0 net6
rlabel metal1 8188 12614 8188 12614 0 net7
rlabel metal1 7498 12614 7498 12614 0 net8
rlabel metal1 2346 11764 2346 11764 0 net9
rlabel metal1 3450 2924 3450 2924 0 next_state\[0\]
rlabel metal1 3450 5780 3450 5780 0 next_state\[1\]
rlabel metal3 1050 10948 1050 10948 0 reset
rlabel metal1 1426 8058 1426 8058 0 spike
rlabel metal2 3634 3876 3634 3876 0 state\[0\]
rlabel metal2 6210 7140 6210 7140 0 state\[1\]
rlabel metal2 6486 1520 6486 1520 0 voltage[0]
rlabel metal2 7130 1520 7130 1520 0 voltage[1]
rlabel metal2 7774 1520 7774 1520 0 voltage[2]
rlabel via2 11914 6171 11914 6171 0 voltage[3]
rlabel metal2 11914 8755 11914 8755 0 voltage[4]
rlabel metal1 6532 12886 6532 12886 0 voltage[5]
rlabel metal1 5842 12954 5842 12954 0 voltage[6]
rlabel metal1 1426 10234 1426 10234 0 voltage[7]
<< properties >>
string FIXED_BBOX 0 0 13499 15643
<< end >>
