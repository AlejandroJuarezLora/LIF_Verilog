magic
tech sky130A
magscale 1 2
timestamp 1727525582
<< nwell >>
rect 1066 2159 12366 13073
<< obsli1 >>
rect 1104 2159 12328 13073
<< obsm1 >>
rect 1104 2128 12328 13104
<< metal2 >>
rect 5814 14843 5870 15643
rect 6458 14843 6514 15643
rect 7102 14843 7158 15643
rect 7746 14843 7802 15643
rect 8390 14843 8446 15643
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
<< obsm2 >>
rect 1306 14787 5758 14843
rect 5926 14787 6402 14843
rect 6570 14787 7046 14843
rect 7214 14787 7690 14843
rect 7858 14787 8334 14843
rect 8502 14787 12034 14843
rect 1306 856 12034 14787
rect 1306 800 5758 856
rect 5926 800 6402 856
rect 6570 800 7046 856
rect 7214 800 7690 856
rect 7858 800 12034 856
<< metal3 >>
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 0 10208 800 10328
rect 12699 9528 13499 9648
rect 12699 8848 13499 8968
rect 0 8168 800 8288
rect 12699 6128 13499 6248
rect 12699 5448 13499 5568
rect 12699 4768 13499 4888
rect 12699 3408 13499 3528
<< obsm3 >>
rect 800 11768 12699 13089
rect 880 11488 12699 11768
rect 800 11088 12699 11488
rect 880 10808 12699 11088
rect 800 10408 12699 10808
rect 880 10128 12699 10408
rect 800 9728 12699 10128
rect 800 9448 12619 9728
rect 800 9048 12699 9448
rect 800 8768 12619 9048
rect 800 8368 12699 8768
rect 880 8088 12699 8368
rect 800 6328 12699 8088
rect 800 6048 12619 6328
rect 800 5648 12699 6048
rect 800 5368 12619 5648
rect 800 4968 12699 5368
rect 800 4688 12619 4968
rect 800 3608 12699 4688
rect 800 3328 12619 3608
rect 800 2143 12699 3328
<< metal4 >>
rect 2347 2128 2667 13104
rect 3007 2128 3327 13104
rect 5153 2128 5473 13104
rect 5813 2128 6133 13104
rect 7959 2128 8279 13104
rect 8619 2128 8939 13104
rect 10765 2128 11085 13104
rect 11425 2128 11745 13104
<< obsm4 >>
rect 4107 8195 4173 11661
<< metal5 >>
rect 1056 12196 12376 12516
rect 1056 11536 12376 11856
rect 1056 9476 12376 9796
rect 1056 8816 12376 9136
rect 1056 6756 12376 7076
rect 1056 6096 12376 6416
rect 1056 4036 12376 4356
rect 1056 3376 12376 3696
<< labels >>
rlabel metal4 s 3007 2128 3327 13104 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5813 2128 6133 13104 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8619 2128 8939 13104 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11425 2128 11745 13104 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4036 12376 4356 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6756 12376 7076 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9476 12376 9796 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12196 12376 12516 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2347 2128 2667 13104 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5153 2128 5473 13104 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7959 2128 8279 13104 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10765 2128 11085 13104 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3376 12376 3696 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6096 12376 6416 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8816 12376 9136 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11536 12376 11856 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 11568 800 11688 6 clk
port 3 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 current[0]
port 4 nsew signal input
rlabel metal3 s 12699 3408 13499 3528 6 current[1]
port 5 nsew signal input
rlabel metal3 s 12699 4768 13499 4888 6 current[2]
port 6 nsew signal input
rlabel metal3 s 12699 5448 13499 5568 6 current[3]
port 7 nsew signal input
rlabel metal3 s 12699 9528 13499 9648 6 current[4]
port 8 nsew signal input
rlabel metal2 s 8390 14843 8446 15643 6 current[5]
port 9 nsew signal input
rlabel metal2 s 7746 14843 7802 15643 6 current[6]
port 10 nsew signal input
rlabel metal2 s 7102 14843 7158 15643 6 current[7]
port 11 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 reset
port 12 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 spike
port 13 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 voltage[0]
port 14 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 voltage[1]
port 15 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 voltage[2]
port 16 nsew signal output
rlabel metal3 s 12699 6128 13499 6248 6 voltage[3]
port 17 nsew signal output
rlabel metal3 s 12699 8848 13499 8968 6 voltage[4]
port 18 nsew signal output
rlabel metal2 s 6458 14843 6514 15643 6 voltage[5]
port 19 nsew signal output
rlabel metal2 s 5814 14843 5870 15643 6 voltage[6]
port 20 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 voltage[7]
port 21 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 13499 15643
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 759940
string GDS_FILE /openlane/designs/LIF/runs/prueba/results/signoff/LIF.magic.gds
string GDS_START 355012
<< end >>

