* NGSPICE file created from LIF.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt LIF VGND VPWR clk current[0] current[1] current[2] current[3] current[4] current[5]
+ current[6] current[7] reset spike voltage[0] voltage[1] voltage[2] voltage[3] voltage[4]
+ voltage[5] voltage[6] voltage[7]
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_200_ _041_ _042_ _044_ _067_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__o211a_1
X_131_ _076_ net6 VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ net16 VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput10 net10 VGND VGND VPWR VPWR spike sky130_fd_sc_hd__buf_2
XFILLER_0_7_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_189_ _103_ _110_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput11 net11 VGND VGND VPWR VPWR voltage[0] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_188_ _093_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput12 net20 VGND VGND VPWR VPWR voltage[1] sky130_fd_sc_hd__buf_2
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_187_ _084_ _086_ _090_ _091_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_18_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_1_1__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_239_ clknet_1_0__leaf_clk _012_ VGND VGND VPWR VPWR next_state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput13 net13 VGND VGND VPWR VPWR voltage[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_186_ _068_ _029_ _031_ _032_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a31oi_1
X_238_ clknet_1_0__leaf_clk _011_ VGND VGND VPWR VPWR next_state\[0\] sky130_fd_sc_hd__dfxtp_1
X_169_ net18 _068_ _114_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR voltage[3] sky130_fd_sc_hd__buf_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_185_ _076_ _067_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_168_ _069_ _101_ _102_ _113_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__a31o_1
X_237_ net9 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR voltage[4] sky130_fd_sc_hd__buf_2
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ _022_ _030_ _109_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a21o_1
X_167_ _109_ _112_ _067_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__o21ai_1
X_236_ net9 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_219_ net8 net7 net6 net5 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput16 net16 VGND VGND VPWR VPWR voltage[5] sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_15_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ _076_ _118_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_3_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_235_ net9 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
X_166_ net18 _111_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_19_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_149_ _070_ _073_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__nor2_1
X_218_ net4 net3 net2 net1 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput17 net17 VGND VGND VPWR VPWR voltage[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_182_ _115_ _027_ _028_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_165_ _104_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__nor2_1
X_234_ net9 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_148_ _084_ _086_ _090_ _091_ _093_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__a311o_2
X_217_ _076_ _075_ _103_ net19 net18 VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__o311a_1
Xoutput18 net18 VGND VGND VPWR VPWR voltage[7] sky130_fd_sc_hd__buf_2
XFILLER_0_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_250_ clknet_1_1__leaf_clk _021_ _010_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_4
X_181_ _026_ _097_ _081_ _094_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__o211a_1
Xfanout20 net12 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_164_ net13 _105_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__and2_1
X_233_ _064_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_216_ _065_ _115_ net23 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a21o_1
X_147_ _081_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ _081_ _094_ _026_ _097_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a211oi_1
X_232_ _064_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_163_ _108_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_215_ _051_ _068_ _055_ _056_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_6_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_146_ _079_ _080_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_129_ net15 VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__buf_1
XFILLER_0_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_231_ _064_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__inv_2
X_162_ net18 _104_ _106_ _107_ state\[1\] VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__o311ai_2
Xinput1 current[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_214_ _107_ net1 _069_ net11 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__o211a_1
X_145_ _080_ _083_ _082_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ _070_ _073_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_161_ state\[0\] VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__inv_2
X_230_ _064_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
Xinput2 current[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_213_ _115_ net1 _109_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__o21ai_1
X_144_ _088_ _086_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nand3_2
X_127_ _071_ _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_160_ net13 _105_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 current[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_212_ net20 _068_ _050_ _054_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__o22a_1
X_143_ net12 net2 _085_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_126_ net19 net7 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 current[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_211_ _065_ _053_ _115_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a21oi_1
X_142_ net11 net1 _087_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_125_ net19 net7 VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 current[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_0_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_210_ _051_ _052_ _088_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_2_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_141_ net20 net2 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__xnor2_1
X_124_ net16 net6 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 current[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_140_ net20 net2 _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ state\[1\] VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 current[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_199_ _035_ _043_ _109_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_122_ _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 current[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_198_ _103_ _110_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_6_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout19 net17 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
Xinput9 reset VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_0_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_197_ _040_ _086_ _090_ state\[1\] VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ _065_ state\[1\] VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__or2_1
X_249_ clknet_1_1__leaf_clk _020_ _009_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 next_state\[1\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_196_ _086_ _090_ _040_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__a21oi_1
X_248_ clknet_1_1__leaf_clk _019_ _008_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
X_179_ _078_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 next_state\[0\] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ _091_ _084_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_247_ clknet_1_1__leaf_clk _018_ _007_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
X_178_ net19 _068_ _025_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 net10 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ _039_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_177_ _115_ _098_ _117_ _024_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_246_ clknet_1_0__leaf_clk _017_ _006_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_229_ _064_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_193_ _075_ _038_ _067_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_245_ clknet_1_0__leaf_clk _016_ _005_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_7_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_176_ _109_ _023_ _067_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_159_ net20 net11 VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__or2_1
X_228_ _064_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_192_ _069_ _094_ _034_ _037_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_244_ clknet_1_0__leaf_clk _015_ _004_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_175_ net19 _022_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_227_ net9 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_158_ net19 _076_ net15 _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_17_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_191_ _118_ _036_ _108_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_243_ clknet_1_0__leaf_clk _014_ _003_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_2
X_174_ _076_ _118_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_226_ _063_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__clkbuf_1
X_157_ net14 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__buf_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_209_ net1 _087_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_17_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_190_ _075_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_242_ clknet_1_0__leaf_clk net21 _002_ VGND VGND VPWR VPWR state\[1\] sky130_fd_sc_hd__dfrtp_2
X_173_ _075_ _103_ _110_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_5_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_156_ _074_ _098_ _100_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__or3_1
X_225_ net21 _065_ _061_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ net11 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__inv_2
X_139_ net13 net3 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__xor2_2
XFILLER_0_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_172_ _116_ _096_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__and2_1
X_241_ clknet_1_0__leaf_clk net22 _001_ VGND VGND VPWR VPWR state\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_224_ _062_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__clkbuf_1
X_155_ _074_ _098_ _100_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__o21ai_1
X_207_ _105_ _049_ _109_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a21oi_1
X_138_ _080_ _082_ _083_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_171_ _078_ _081_ _094_ _097_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__a31o_1
X_240_ clknet_1_1__leaf_clk _013_ _000_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_223_ net22 _069_ _061_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__mux2_1
X_154_ _071_ _099_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__xnor2_1
X_206_ net20 net11 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2_1
X_137_ net13 net3 VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_170_ state\[1\] VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_153_ net18 net8 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__xor2_1
X_222_ _107_ state\[1\] _057_ _060_ _000_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_9_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_205_ net13 _107_ _069_ _047_ _048_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a311o_1
X_136_ net14 net4 VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_119_ state\[0\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_152_ _078_ _081_ _094_ _096_ _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__a311oi_2
X_221_ net9 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_204_ _065_ _110_ _106_ _115_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and4bb_1
X_135_ _079_ _080_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_220_ _066_ _058_ _059_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__or3_1
X_151_ _075_ net5 _070_ _077_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_203_ _065_ _069_ _090_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__and4_1
X_134_ net14 net4 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_150_ _074_ _095_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ _086_ _089_ _088_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a21o_1
X_133_ net15 net5 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_201_ _103_ _068_ _045_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__o21ba_1
X_132_ _075_ net5 _070_ _077_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_16_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

